DirectoryBRAM.bsv