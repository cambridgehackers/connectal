/* Copyright (c) 2014 Quanta Research Cambridge, Inc
 *
 * Permission is hereby granted, free of charge, to any person obtaining a
 * copy of this software and associated documentation files (the "Software"),
 * to deal in the Software without restriction, including without limitation
 * the rights to use, copy, modify, merge, publish, distribute, sublicense,
 * and/or sell copies of the Software, and to permit persons to whom the
 * Software is furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included
 * in all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
 * OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
 * FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
 * DEALINGS IN THE SOFTWARE.
 */
// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;
import BRAM::*;
import DefaultValue::*;
import Connectable::*;

// connectal libraries
import Leds::*;
import CtrlMux::*;
import Portal::*;
import ConnectalMemory::*;
import MemTypes::*;
import MemServer::*;
import MemServerInternal::*;
import MMU::*;
import MemreadEngine::*;
import MemwriteEngine::*;
import HostInterface::*;

// generated by tool
import MMURequest::*;
import StrstrRequest::*;
import MemServerIndication::*;
import MMUIndication::*;
import StrstrIndication::*;


import Strstr::*;
// import AuroraCommon::*;
// import FlashTop::*;
// import FlashRequest::*;
// import FlashIndication::*;

typedef enum {
   FlashIndication, 
   FlashRequest, 

   HostMemServerIndication, 
   HostMemServerRequest, 
   
   FlashMemServerIndication, 
   FlashMemServerRequest, 
	      
   HostMMURequest, 
   HostMMUIndication, 

   FlashMMURequest, 
   FlashMMUIndication,

   AlgoIndication, 
   AlgoRequest 

} IfcNames deriving (Eq,Bits);

// interface Top_Pins;
// 	interface Aurora_Pins#(4) aurora_fmc1;
// 	interface Aurora_Clock_Pins aurora_clk_fmc1;
// endinterface

typedef 128 FlashDataWidth;
typedef 30  FlashAddrWidth;

//module mkConnectalTop#(HostType host) (StdConnectalDmaTop#(PhysAddrWidth));
module mkConnectalTop(StdConnectalDmaTop#(PhysAddrWidth));
   
   // Clock clk250 = host.doubleClock;
   // Reset rst250 = host.doubleReset;
	
   // strstr algo
   StrstrIndicationProxy strstrIndicationProxy <- mkStrstrIndicationProxy(AlgoIndication);
   Strstr#(128,64) strstr <- mkStrstr(strstrIndicationProxy.ifc);
   StrstrRequestWrapper strstrRequestWrapper <- mkStrstrRequestWrapper(AlgoRequest,strstr.request);
   
   // host mmu
   MMUIndicationProxy hostMMUIndicationProxy <- mkMMUIndicationProxy(HostMMUIndication);
   MMU#(PhysAddrWidth) hostMMU <- mkMMU(1, True, hostMMUIndicationProxy.ifc);
   MMURequestWrapper hostMMURequestWrapper <- mkMMURequestWrapper(HostMMURequest, hostMMU.request);
   
   // flash mmu
   MMUIndicationProxy flashMMUIndicationProxy <- mkMMUIndicationProxy(FlashMMUIndication);
   MMU#(FlashAddrWidth) flashMMU <- mkMMU(0, False, flashMMUIndicationProxy.ifc);
   MMURequestWrapper flashMMURequestWrapper <- mkMMURequestWrapper(FlashMMURequest, flashMMU.request);

   // flash top
   // FlashIndicationProxy flashIndicationProxy <- mkFlashIndicationProxy(FlashIndication);
   // FlashTop flashtop <- mkFlashTop(flashIndicationProxy.ifc, clk250, rst250);
   // FlashRequestWrapper flashRequestWrapper <- mkFlashRequestWrapper(FlashRequest,flashtop.request);
   
   // host memory server
   MemServerIndicationProxy hostMemServerIndicationProxy <- mkMemServerIndicationProxy(HostMemServerIndication);
   let rcs = cons(strstr.config_read_client,nil);//cons(flashtop.hostMemReadClient,nil));
   //let wcs = cons(flashtop.hostMemWriteClient,nil);
   let mmus = cons(hostMMU,nil);
   //MemServer#(PhysAddrWidth,64,1) hostMemServer <- mkMemServerRW(hostMemServerIndicationProxy.ifc, rcs, wcs, mmus);
   MemServer#(PhysAddrWidth,64,1) hostMemServer <- mkMemServerR(hostMemServerIndicationProxy.ifc, rcs, mmus);

   // flash memory read server
   MemServerIndicationProxy flashMemServerIndicationProxy <- mkMemServerIndicationProxy(FlashMemServerIndication);
   MemServer#(FlashAddrWidth,FlashDataWidth,1) flashMemServer <- mkMemServerR(flashMemServerIndicationProxy.ifc, cons(strstr.haystack_read_client,nil),  cons(flashMMU,nil));
   //mkConnection(flashMemServer.masters[0], flashtop.memSlave);
   
   
   Vector#(10,StdPortal) portals;

   portals[0] = strstrRequestWrapper.portalIfc;
   portals[1] = strstrIndicationProxy.portalIfc; 

   portals[2] = hostMMURequestWrapper.portalIfc;
   portals[3] = hostMMUIndicationProxy.portalIfc;
   
   portals[4] = flashMMURequestWrapper.portalIfc;
   portals[5] = flashMMUIndicationProxy.portalIfc; 
   
   portals[6] = ?; //flashRequestWrapper.portalIfc;
   portals[7] = ?; //flashIndicationProxy.portalIfc;
   
   portals[8] = hostMemServerIndicationProxy.portalIfc;
   portals[9] = flashMemServerIndicationProxy.portalIfc;
   
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = hostMemServer.masters;
   interface leds = default_leds;
      
endmodule : mkConnectalTop


