// bsv libraries
import Vector::*;
import FIFO::*;
import Connectable::*;
import Portal::*;
import CtrlMux::*;
import Leds::*;
import MemTypes::*;
import MMU::*;
import MemServer::*;
import MemPortal::*;

// generated by tool
import EchoIndication::*;
import EchoRequest::*;
import Swallow::*;

import DmaDebugRequest::*;
import MMUConfigRequest::*;
import DmaDebugIndication::*;
import MMUConfigIndication::*;
import MMUConfigIndication::*;
import SharedMemoryPortalConfig::*;

// defined by user
import Echo::*;
import SwallowIF::*;

typedef enum {EchoIndication, EchoRequest, Swallow, SS_EchoRequest, SS_EchoIndication,
MMUConfigRequest, MMUConfigIndication, DmaDebugIndication, DmaDebugRequest, ConfigWrapper} IfcNames deriving (Eq,Bits);

module mkConnectalTop(StdConnectalDmaTop#(PhysAddrWidth));

   // instantiate user portals
   EchoIndicationProxy echoIndicationProxy <- mkEchoIndicationProxy(EchoIndication);
   EchoRequestInternal echoRequestInternal <- mkEchoRequestInternal(echoIndicationProxy.ifc);
   EchoRequestWrapperPortal echoRequestWrapper <- mkEchoRequestWrapperPortal(EchoRequest,echoRequestInternal.ifc);
   
   Swallow swallow <- mkSwallow();
   SwallowWrapper swallowWrapper <- mkSwallowWrapper(Swallow, swallow);
   
   SharedMemoryPortal#(64) echoRequestSharedMemoryPortal <- mkSharedMemoryPortal(echoRequestWrapper.portalIfc);
   SharedMemoryPortalConfigWrapper configWrapper <- mkSharedMemoryPortalConfigWrapper(ConfigWrapper, echoRequestSharedMemoryPortal.cfg);

   let readClients = cons(echoRequestSharedMemoryPortal.readClient, nil);
   let writeClients = cons(echoRequestSharedMemoryPortal.writeClient, nil);

   MMUConfigIndicationProxy mmuConfigIndicationProxy <- mkMMUConfigIndicationProxy(MMUConfigIndication);
   MMU#(PhysAddrWidth) mmu <- mkMMU(0, True, mmuConfigIndicationProxy.ifc);
   MMUConfigRequestWrapper mmuConfigRequestWrapper <- mkMMUConfigRequestWrapper(MMUConfigRequest, mmu.request);

   DmaDebugIndicationProxy dmaDebugIndicationProxy <- mkDmaDebugIndicationProxy(DmaDebugIndication);
   MemServer#(PhysAddrWidth,64,1) dma <- mkMemServerRW(dmaDebugIndicationProxy.ifc, readClients, writeClients, cons(mmu,nil));
   DmaDebugRequestWrapper dmaDebugRequestWrapper <- mkDmaDebugRequestWrapper(DmaDebugRequest, dma.request);

   Vector#(7,StdPortal) portals;
   portals[0] = swallowWrapper.portalIfc;
   portals[1] = echoIndicationProxy.portalIfc;
   portals[2] = dmaDebugIndicationProxy.portalIfc; 
   portals[3] = dmaDebugRequestWrapper.portalIfc;
   portals[4] = mmuConfigRequestWrapper.portalIfc;
   portals[5] = mmuConfigIndicationProxy.portalIfc;
   portals[6] = configWrapper.portalIfc;
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = echoRequestInternal.leds;
   interface Empty pins;
   endinterface

endmodule : mkConnectalTop
