// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import Directory::*;
import CtrlMux::*;
import Portal::*;
import PortalMemory::*;
import MemTypes::*;
import DmaUtils::*;
import MemServer::*;

// generated by tool
import Memread2RequestWrapper::*;
import DmaConfigWrapper::*;
import Memread2IndicationProxy::*;
import DmaIndicationProxy::*;

// defined by user
import Memread2::*;

typedef enum {Memread2Indication, Memread2Request, DmaIndication, DmaConfig} IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalDmaTop#(addrWidth)) provisos (
    Add#(addrWidth, a__, 52),
    Add#(b__, addrWidth, 64),
    Add#(c__, 12, addrWidth),
    Add#(addrWidth, d__, 44),
    Add#(e__, addrWidth, 40),
    Add#(f__, c__, 40));

   DmaIndicationProxy dmaIndicationProxy <- mkDmaIndicationProxy(DmaIndication);

   Memread2IndicationProxy memreadIndicationProxy <- mkMemread2IndicationProxy(Memread2Indication);
   Memread2 memread <- mkMemread2(memreadIndicationProxy.ifc);
   Memread2RequestWrapper memreadRequestWrapper <- mkMemread2RequestWrapper(Memread2Request,memread.request);

   Vector#(2, ObjectReadClient#(64)) clients;
   Vector#(2, DmaReadBuffer#(64, 16)) readBuffers <- replicateM(mkDmaReadBuffer);
   mkConnection(memread.dmaClient, readBuffers[0].dmaServer);
   mkConnection(memread.dmaClient2, readBuffers[1].dmaServer);
   clients = cons(readBuffers[0].dmaClient, cons(readBuffers[1].dmaClient, nil));
   MemServer#(addrWidth,64,1) dma <- mkMemServerR(dmaIndicationProxy.ifc, clients);

   DmaConfigWrapper dmaRequestWrapper <- mkDmaConfigWrapper(DmaConfig,dma.request);

   Vector#(4,StdPortal) portals;
   portals[0] = memreadRequestWrapper.portalIfc;
   portals[1] = memreadIndicationProxy.portalIfc; 
   portals[2] = dmaRequestWrapper.portalIfc;
   portals[3] = dmaIndicationProxy.portalIfc; 
   
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = ?;
endmodule : mkPortalTop
