// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import AxiMasterSlave::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import PortalMemory::*;
import Dma::*;
import AxiDma::*;
import Leds::*;
import DmaUtils::*;
import HDMI::*;

// generated by tool
import DmaConfigWrapper::*;
import DmaIndicationProxy::*;
import HdmiControlRequestWrapper::*;
import HdmiInternalIndicationProxy::*;
import HdmiInternalRequestWrapper::*;

// defined by user
import HdmiDisplay::*;

typedef enum {HdmiControlRequest, HdmiInternalRequest, HdmiInternalIndication, DmaConfig, DmaIndication} IfcNames deriving (Eq,Bits);

module mkPortalTop#(Clock clk1)(PortalTop#(addrWidth,64,HDMI))
   provisos(Add#(addrWidth, a__, 52),
	    Add#(b__, addrWidth, 64),
	    Add#(c__, 12, addrWidth),
	    Add#(addrWidth, d__, 44),
	    Add#(e__, c__, DmaOffsetSize),
	    Add#(f__, addrWidth, 40));

   HdmiInternalIndicationProxy hdmiInternalIndicationProxy <- mkHdmiInternalIndicationProxy(HdmiInternalIndication);
   HdmiDisplay hdmiDisplay <- mkHdmiDisplay(clk1, hdmiInternalIndicationProxy.ifc);
   HdmiControlRequestWrapper hdmiControlRequestWrapper <- mkHdmiControlRequestWrapper(HdmiControlRequest,hdmiDisplay.controlRequest);
   HdmiInternalRequestWrapper hdmiInternalRequestWrapper <- mkHdmiInternalRequestWrapper(HdmiInternalRequest,hdmiDisplay.internalRequest);

   DmaIndicationProxy dmaIndicationProxy <- mkDmaIndicationProxy(DmaIndication);
   Vector#(1,  DmaReadClient#(64))   readClients = cons(hdmiDisplay.dmaClient, nil);
   Integer               numRequests = 8;
   AxiDmaServer#(addrWidth, 64)   dma <- mkAxiDmaServer(dmaIndicationProxy.ifc, numRequests, readClients, nil);
   DmaConfigWrapper dmaRequestWrapper <- mkDmaConfigWrapper(DmaConfig,dma.request);

   Vector#(5,StdPortal) portals;
   portals[0] = hdmiControlRequestWrapper.portalIfc;
   portals[1] = hdmiInternalRequestWrapper.portalIfc;
   portals[2] = hdmiInternalIndicationProxy.portalIfc; 
   portals[3] = dmaRequestWrapper.portalIfc;
   portals[4] = dmaIndicationProxy.portalIfc; 
   
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkAxiSlaveMux(dir,portals);
   let interrupt_mux <- mkInterruptMux(portals);
   
   interface interrupt = interrupt_mux;
   interface ctrl = ctrl_mux;
   interface m_axi = dma.m_axi;
   interface leds = default_leds;
      
endmodule : mkPortalTop
