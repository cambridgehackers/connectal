// bsv libraries
import Vector::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import Portal::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import AxiMasterSlave::*;

// generated by tool
import ImageCaptureIndicationProxy::*;
import ImageCaptureRequestWrapper::*;

// defined by user
import ImageCapture::*;

typedef enum {ImageCaptureIndication, ImageCaptureRequest} IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalTop#(addrWidth));

   // instantiate user portals
   ImageCaptureIndicationProxy captureIndicationProxy <- mkImageCaptureIndicationProxy(ImageCaptureIndication);
   ImageCaptureRequestInternal captureRequestInternal <- mkImageCaptureRequestInternal(captureIndicationProxy.ifc);
   ImageCaptureRequestWrapper captureRequestWrapper <- mkImageCaptureRequestWrapper(ImageCaptureRequest,captureRequestInternal.ifc);
   
   ImageCaptureRequest capture <- mkImageCaptureRequest();
   ImageCaptureWrapper captureWrapper <- mkImageCaptureWrapper(ImageCapture, capture);
   
   Vector#(3,StdPortal) portals;
   portals[0] = captureIndicationProxy.portalIfc;
   portals[1] = captureRequestWrapper.portalIfc; 
   portals[2] = captureWrapper.portalIfc; 
   let interrupt_mux <- mkInterruptMux(portals);
   
   // instantiate system directory
   Directory dir <- mkDirectoryDbg(portals,interrupt_mux);
   Vector#(1,StdPortal) directories;
   directories[0] = dir.portalIfc;
   
   // when constructing the ctrl mux, directories must be the first argument
   let ctrl_mux <- mkAxiSlaveMux(directories,portals);
   
   interface interrupt = interrupt_mux;
   interface ctrl = ctrl_mux;
   interface m_axi = null_axi_master;
   interface leds = captureRequestInternal.leds;

endmodule : mkPortalTop
