// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;
import BRAM::*;
import DefaultValue::*;
import Connectable::*;

// portz libraries
import Leds::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import PortalMemory::*;
import MemTypes::*;
import MemServer::*;
import MemServerInternal::*;
import SGList::*;


// generated by tool
import NandSimRequestWrapper::*;
import DmaConfigWrapper::*;
import StrstrRequestWrapper::*;

import NandSimIndicationProxy::*;
import DmaIndicationProxy::*;
import StrstrIndicationProxy::*;

// defined by user
import NandSim::*;
import NandSimNames::*;
import Strstr::*;

`ifdef BSIM
`ifndef PCIE
import "BDPI" function ActionValue#(Bit#(32)) pareff_init(Bit#(32) id, Bit#(32) handle, Bit#(32) size);
`endif
`endif

module mkPortalTop(StdPortalDmaTop#(PhysAddrWidth));
   
   NandSimIndicationProxy nandSimIndicationProxy <- mkNandSimIndicationProxy(NandSimIndication);
   NandSim nandSim <- mkNandSim(nandSimIndicationProxy.ifc);
   NandSimRequestWrapper nandSimRequestWrapper <- mkNandSimRequestWrapper(NandSimRequest,nandSim.request);
   
   StrstrIndicationProxy strstrIndicationProxy <- mkStrstrIndicationProxy(AlgoIndication);
   Strstr#(1,64) strstr <- mkStrstr(strstrIndicationProxy.ifc);
   StrstrRequestWrapper strstrRequestWrapper <- mkStrstrRequestWrapper(AlgoRequest,strstr.request);
   
   DmaIndicationProxy dmaIndicationProxy <- mkDmaIndicationProxy(DmaIndication);
   let rcs = cons(strstr.config_read_client,cons(nandSim.readClient, nil));
   SGListMMU#(PhysAddrWidth) sgl0 <- mkSGListMMU(0, True, dmaIndicationProxy.ifc);
   MemServer#(PhysAddrWidth,64,1) dma <- mkConfigMemServerRW(dmaIndicationProxy.ifc, rcs, cons(nandSim.writeClient, nil), sgl0);
   DmaConfigWrapper dmaRequestWrapper <- mkDmaConfigWrapper(DmaConfig, dma.request);

   DmaIndicationProxy nandsimDmaIndicationProxy <- mkDmaIndicationProxy(NandsimDmaIndication);   
   SGListMMU#(PhysAddrWidth) sgl1 <- mkSGListMMU(1, False, nandsimDmaIndicationProxy.ifc);
   MemServer#(PhysAddrWidth,64,1) nandsimDma <- mkConfigMemServerR(nandsimDmaIndicationProxy.ifc, cons(strstr.haystack_read_client,nil), sgl1);
   DmaConfigWrapper nandsimDmaRequestWrapper <- mkDmaConfigWrapper(NandsimDmaConfig, nandsimDma.request);
   mkConnection(nandsimDma.masters[0], nandSim.memSlave);
   
   
   Vector#(8,StdPortal) portals;
   portals[0] = nandSimRequestWrapper.portalIfc;
   portals[1] = nandSimIndicationProxy.portalIfc; 
   portals[2] = dmaRequestWrapper.portalIfc;
   portals[3] = dmaIndicationProxy.portalIfc; 
   portals[4] = strstrRequestWrapper.portalIfc;
   portals[5] = strstrIndicationProxy.portalIfc; 
   portals[6] = nandsimDmaRequestWrapper.portalIfc;
   portals[7] = nandsimDmaIndicationProxy.portalIfc; 
   
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;
      
endmodule : mkPortalTop
