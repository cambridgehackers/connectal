// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;


// portz libraries
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import PortalMemory::*;
import MemServer::*;
import Dma::*;
import DmaUtils::*;

// generated by tool
import MempokeRequestWrapper::*;
import DmaConfigWrapper::*;
import MempokeIndicationProxy::*;
import DmaIndicationProxy::*;

// defined by user
import Mempoke::*;

typedef enum {MempokeIndication, MempokeRequest, DmaIndication, DmaConfig} IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalDmaTop#(addrWidth)) 

   provisos(Add#(addrWidth, a__, 52),
	    Add#(b__, addrWidth, 64),
	    Add#(c__, 12, addrWidth),
	    Add#(addrWidth, d__, 44),
	    Add#(e__, c__, 40),
	    Add#(f__, addrWidth, 40));

   DmaIndicationProxy dmaIndicationProxy <- mkDmaIndicationProxy(DmaIndication);
   DmaWriteBuffer#(64,16) dma_stream_write_chan <- mkDmaWriteBuffer();
   DmaReadBuffer#(64,16) dma_stream_read_chan <- mkDmaReadBuffer();

   Vector#(1, ObjectReadClient#(64))   readClients = newVector();
   Vector#(1, ObjectWriteClient#(64)) writeClients = newVector();
   writeClients[0] = dma_stream_write_chan.dmaClient;
   readClients[0]  = dma_stream_read_chan.dmaClient;
   MemServer#(addrWidth,64,1)   dma <- mkMemServer(dmaIndicationProxy.ifc, readClients, writeClients);
   DmaConfigWrapper dmaRequestWrapper <- mkDmaConfigWrapper(DmaConfig,dma.request);

   
   MempokeIndicationProxy mempokeIndicationProxy <- mkMempokeIndicationProxy(MempokeIndication);
   MempokeRequest mempokeRequest <- mkMempokeRequest(mempokeIndicationProxy.ifc, dma_stream_write_chan.dmaServer, dma_stream_read_chan.dmaServer);
   MempokeRequestWrapper mempokeRequestWrapper <- mkMempokeRequestWrapper(MempokeRequest,mempokeRequest);

   Vector#(4,StdPortal) portals;
   portals[0] = mempokeRequestWrapper.portalIfc;
   portals[1] = mempokeIndicationProxy.portalIfc; 
   portals[2] = dmaRequestWrapper.portalIfc;
   portals[3] = dmaIndicationProxy.portalIfc; 
   
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;
endmodule
