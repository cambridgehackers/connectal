/* Copyright (c) 2014 Quanta Research Cambridge, Inc
 *
 * Permission is hereby granted, free of charge, to any person obtaining a
 * copy of this software and associated documentation files (the "Software"),
 * to deal in the Software without restriction, including without limitation
 * the rights to use, copy, modify, merge, publish, distribute, sublicense,
 * and/or sell copies of the Software, and to permit persons to whom the
 * Software is furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included
 * in all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
 * OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
 * FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
 * DEALINGS IN THE SOFTWARE.
 */
// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;
import BRAM::*;
import DefaultValue::*;
import Connectable::*;

// portz libraries
import Leds::*;
import CtrlMux::*;
import Portal::*;
import ConnectalMemory::*;
import MemTypes::*;
import MemServer::*;
import MemServerInternal::*;
import MMU::*;


// generated by tool
import NandSimRequest::*;
import MMURequest::*;
import StrstrRequest::*;

import NandSimIndication::*;
import MemServerIndication::*;
import MMUIndication::*;
import StrstrIndication::*;

// defined by user
import NandSim::*;
import NandSimNames::*;
import Strstr::*;

typedef HaystackReadClients NandSimSlaves;

module mkConnectalTop(StdConnectalDmaTop#(PhysAddrWidth));
   
   // nandsim 
   NandSimIndicationProxy nandSimIndicationProxy <- mkNandSimIndicationProxy(NandSimIndication);
   NandSim#(NandSimSlaves) nandSim <- mkNandSim(nandSimIndicationProxy.ifc);
   NandSimRequestWrapper nandSimRequestWrapper <- mkNandSimRequestWrapper(NandSimRequest,nandSim.request);
   
   // strstr algo
   StrstrIndicationProxy strstrIndicationProxy <- mkStrstrIndicationProxy(AlgoIndication);
   Strstr#(64) strstr <- mkStrstr(strstrIndicationProxy.ifc);
   StrstrRequestWrapper strstrRequestWrapper <- mkStrstrRequestWrapper(AlgoRequest,strstr.request);
   
   // backing store mmu
   MMUIndicationProxy backingStoreMMUIndicationProxy <- mkMMUIndicationProxy(BackingStoreMMUIndication);
   MMU#(PhysAddrWidth) backingStoreMMU <- mkMMU(0, True, backingStoreMMUIndicationProxy.ifc);
   MMURequestWrapper backingStoreMMURequestWrapper <- mkMMURequestWrapper(BackingStoreMMURequest, backingStoreMMU.request);

   // algo mmu
   MMUIndicationProxy algoMMUIndicationProxy <- mkMMUIndicationProxy(AlgoMMUIndication);
   MMU#(PhysAddrWidth) algoMMU <- mkMMU(1, True, algoMMUIndicationProxy.ifc);
   MMURequestWrapper algoMMURequestWrapper <- mkMMURequestWrapper(AlgoMMURequest, algoMMU.request);
      
   // host memory dma server
   MemServerIndicationProxy hostMemServerIndicationProxy <- mkMemServerIndicationProxy(HostMemServerIndication);
   let rcs = cons(strstr.config_read_client,cons(nandSim.readClient, nil));
   MemServer#(PhysAddrWidth,64,1) hostDma <- mkMemServerRW(hostMemServerIndicationProxy.ifc,rcs, cons(nandSim.writeClient, nil), cons(backingStoreMMU,cons(algoMMU,nil)));

   // nandsim mmu0
   MMUIndicationProxy nandsimMMU0IndicationProxy <- mkMMUIndicationProxy(NandsimMMU0Indication);
   MMU#(PhysAddrWidth) nandsimMMU0 <- mkMMU(0, False, nandsimMMU0IndicationProxy.ifc);
   MMURequestWrapper nandsimMMU0RequestWrapper <- mkMMURequestWrapper(NandsimMMU0Request, nandsimMMU0.request);
   
   // nandsim memory dma0 server
   MemServerIndicationProxy nandsimMemServer0IndicationProxy <- mkMemServerIndicationProxy(NandsimMemServer0Indication);   
   MemServer#(PhysAddrWidth,64,1) nandsimDma0 <- mkMemServerR(nandsimMemServer0IndicationProxy.ifc, cons(strstr.haystack_read_clients[0],nil), cons(nandsimMMU0,nil));
   mkConnection(nandsimDma0.masters[0], nandSim.memSlaves[0]);
   
   // nandsim mmu1
   MMUIndicationProxy nandsimMMU1IndicationProxy <- mkMMUIndicationProxy(NandsimMMU1Indication);
   MMU#(PhysAddrWidth) nandsimMMU1 <- mkMMU(0, False, nandsimMMU1IndicationProxy.ifc);
   MMURequestWrapper nandsimMMU1RequestWrapper <- mkMMURequestWrapper(NandsimMMU1Request, nandsimMMU1.request);
   
   // nandsim memory dma1 server
   MemServerIndicationProxy nandsimMemServer1IndicationProxy <- mkMemServerIndicationProxy(NandsimMemServer1Indication);   
   MemServer#(PhysAddrWidth,64,1) nandsimDma1 <- mkMemServerR(nandsimMemServer1IndicationProxy.ifc, cons(strstr.haystack_read_clients[1],nil), cons(nandsimMMU1,nil));
   mkConnection(nandsimDma1.masters[0], nandSim.memSlaves[1]);
   
   Vector#(15,StdPortal) portals;

   portals[0] = nandSimRequestWrapper.portalIfc;
   portals[1] = nandSimIndicationProxy.portalIfc; 

   portals[2] = strstrRequestWrapper.portalIfc;
   portals[3] = strstrIndicationProxy.portalIfc; 
   
   portals[4] = backingStoreMMURequestWrapper.portalIfc;
   portals[5] = backingStoreMMUIndicationProxy.portalIfc;

   portals[6] = algoMMURequestWrapper.portalIfc;
   portals[7] = algoMMUIndicationProxy.portalIfc;
   
   portals[8] = nandsimMMU0RequestWrapper.portalIfc;
   portals[9] = nandsimMMU0IndicationProxy.portalIfc;

   portals[10] = nandsimMMU1RequestWrapper.portalIfc;
   portals[11] = nandsimMMU1IndicationProxy.portalIfc;

   portals[12] = hostMemServerIndicationProxy.portalIfc;
   portals[13] = nandsimMemServer0IndicationProxy.portalIfc;
   portals[14] = nandsimMemServer1IndicationProxy.portalIfc;

   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = hostDma.masters;
   interface leds = default_leds;
      
endmodule : mkConnectalTop
