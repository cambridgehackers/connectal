`define ConnectalVersion 15.10.3
`define NumberOfMasters 1
`define PinType Empty
`define PinTypeInclude Misc
`define NumberOfUserTiles 1
`define SlaveDataBusWidth 32
`define SlaveControlAddrWidth 5
`define BurstLenSize 8
`define project_dir $(DTOP)
`define MainClockPeriod 20
`define DerivedClockPeriod 10.000000
`define BsimHostInterface 
`define PhysAddrWidth 40
`define SIMULATION 
`define BOARD_bluesim 
