// Copyright (c) 2015 Quanta Research Cambridge, Inc.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.


typedef struct {
   t1 tpl_1;
   t2 tpl_2;
   } Tuple2#(type t1, type t2);

typedef struct {
   t1 tpl_1;
   t2 tpl_2;
   t3 tpl_3;
   } Tuple3#(type t1, type t2, type t3);

typedef struct {
   t1 tpl_1;
   t2 tpl_2;
   t3 tpl_3;
   t4 tpl_4;
   } Tuple4#(type t1, type t2, type t3, type t4);

typedef struct {
   t1 tpl_1;
   t2 tpl_2;
   t3 tpl_3;
   t4 tpl_4;
   t5 tpl_5;
   } Tuple5#(type t1, type t2, type t3, type t4, type t5);

