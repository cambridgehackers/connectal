module l_class_OC_Fifo (
    input CLK,
    input nRST);

   reg[31:0]  (**) ( VERILOG_int, ...);
  always @( posedge CLK) begin
    if (!nRST) begin
    end
    else begin
    end; // nRST
  end; // always @ (posedge CLK)
endmodule 

