// bsv libraries
import Vector::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import CtrlMux::*;
import Portal::*;
import Leds::*;
import MemTypes::*;
import MMU::*;
import MemServer::*;
import MemPortal::*;

// generated by tool
import Simple::*;

import MMUConfigRequest::*;
import MMUConfigIndication::*;
import MMUConfigIndication::*;
import SharedMemoryPortalConfig::*;
import DmaDebugIndication::*;

// defined by user
import SimpleIF::*;

typedef enum {SimpleIndication, SimpleRequest,
	      MMUConfigRequest, MMUConfigIndication, DmaDebugIndication, ConfigWrapper} IfcNames deriving (Eq,Bits);

module mkConnectalTop(StdConnectalDmaTop#(PhysAddrWidth));

   // instantiate user portals
   SimpleProxy simpleIndicationProxy <- mkSimpleProxy(SimpleIndication);
   Simple simpleRequest <- mkSimple(simpleIndicationProxy.ifc);
   SimpleWrapperPortal simpleRequestWrapper <- mkSimpleWrapperPortal(SimpleRequest,simpleRequest);
   
   SharedMemoryPortal#(64) echoRequestSharedMemoryPortal <- mkSharedMemoryPortal(simpleRequestWrapper.portalIfc);
   SharedMemoryPortalConfigWrapper configWrapper <- mkSharedMemoryPortalConfigWrapper(ConfigWrapper, echoRequestSharedMemoryPortal.cfg);

   let readClients = cons(echoRequestSharedMemoryPortal.readClient, nil);
   let writeClients = cons(echoRequestSharedMemoryPortal.writeClient, nil);

   DmaDebugIndicationProxy dmaDebugIndicationProxy <- mkDmaDebugIndicationProxy(DmaDebugIndication);
   MMUConfigIndicationProxy mmuConfigIndicationProxy <- mkMMUConfigIndicationProxy(MMUConfigIndication);
   MMU#(PhysAddrWidth) mmu <- mkMMU(0, True, mmuConfigIndicationProxy.ifc);
   MMUConfigRequestWrapper mmuConfigRequestWrapper <- mkMMUConfigRequestWrapper(MMUConfigRequest, mmu.request);
   MemServer#(PhysAddrWidth,64,1) dma <- mkMemServerRW(mmuConfigIndicationProxy.ifc, dmaDebugIndicationProxy.ifc, readClients, writeClients, cons(mmu,nil));

   Vector#(5,StdPortal) portals;
   portals[0] = simpleIndicationProxy.portalIfc;
   portals[1] = mmuConfigRequestWrapper.portalIfc;
   portals[2] = mmuConfigIndicationProxy.portalIfc;
   portals[3] = configWrapper.portalIfc;
   portals[4] = dmaDebugIndicationProxy.portalIfc;
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;

endmodule : mkConnectalTop


