// bsv libraries
import Vector::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import CtrlMux::*;
import Portal::*;
import Leds::*;
import MemTypes::*;
import MemPortal::*;

// generated by tool
import MifoTestIndication::*;
import MifoTestRequest::*;

// defined by user
import MifoTest::*;

typedef enum {MifoTestIndication, MifoTestRequest} IfcNames deriving (Eq,Bits);

module mkConnectalTop(StdConnectalTop#(PhysAddrWidth));

   // instantiate user portals
   MifoTestIndicationProxy mifoIndicationProxy <- mkMifoTestIndicationProxy(MifoTestIndication);
   MifoTestRequest mifoRequest <- mkMifoTestRequest(mifoIndicationProxy.ifc);
   MifoTestRequestWrapper mifoRequestWrapper <- mkMifoTestRequestWrapper(MifoTestRequest,mifoRequest);
   
   Vector#(2,StdPortal) portals;
   portals[0] = mifoRequestWrapper.portalIfc;
   portals[1] = mifoIndicationProxy.portalIfc;
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = nil;
   interface leds = default_leds;

endmodule : mkConnectalTop


