
typedef enum {IfcNames_MemwriteIndicationH2S, IfcNames_MemwriteRequestS2H} TileNames deriving (Eq,Bits);
