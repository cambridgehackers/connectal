// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;
import BRAM::*;
import DefaultValue::*;
import Connectable::*;

// portz libraries
import Leds::*;
import CtrlMux::*;
import Portal::*;
import ConnectalMemory::*;
import MemTypes::*;
import MemServer::*;
import MemServerInternal::*;
import MMU::*;


// generated by tool
import NandSimRequest::*;
import MMUConfigRequest::*;
import StrstrRequest::*;

import NandSimIndication::*;
import DmaDebugIndication::*;
import MMUConfigIndication::*;
import StrstrIndication::*;

// defined by user
import NandSim::*;
import NandSimNames::*;
import Strstr::*;

typedef HaystackReadClients NandSimSlaves;

module mkConnectalTop(StdConnectalDmaTop#(PhysAddrWidth));
   
   // nandsim 
   NandSimIndicationProxy nandSimIndicationProxy <- mkNandSimIndicationProxy(NandSimIndication);
   NandSim#(NandSimSlaves) nandSim <- mkNandSim(nandSimIndicationProxy.ifc);
   NandSimRequestWrapper nandSimRequestWrapper <- mkNandSimRequestWrapper(NandSimRequest,nandSim.request);
   
   // strstr algo
   StrstrIndicationProxy strstrIndicationProxy <- mkStrstrIndicationProxy(AlgoIndication);
   Strstr#(64) strstr <- mkStrstr(strstrIndicationProxy.ifc);
   StrstrRequestWrapper strstrRequestWrapper <- mkStrstrRequestWrapper(AlgoRequest,strstr.request);
   
   // backing store mmu
   MMUConfigIndicationProxy backingStoreMMUConfigIndicationProxy <- mkMMUConfigIndicationProxy(BackingStoreMMUConfigIndication);
   MMU#(PhysAddrWidth) backingStoreMMU <- mkMMU(0, True, backingStoreMMUConfigIndicationProxy.ifc);
   MMUConfigRequestWrapper backingStoreMMUConfigRequestWrapper <- mkMMUConfigRequestWrapper(BackingStoreMMUConfigRequest, backingStoreMMU.request);

   // algo mmu
   MMUConfigIndicationProxy algoMMUConfigIndicationProxy <- mkMMUConfigIndicationProxy(AlgoMMUConfigIndication);
   MMU#(PhysAddrWidth) algoMMU <- mkMMU(1, True, algoMMUConfigIndicationProxy.ifc);
   MMUConfigRequestWrapper algoMMUConfigRequestWrapper <- mkMMUConfigRequestWrapper(AlgoMMUConfigRequest, algoMMU.request);
      
   // host memory dma server
   DmaDebugIndicationProxy hostDmaDebugIndicationProxy <- mkDmaDebugIndicationProxy(HostDmaDebugIndication);
   let rcs = cons(strstr.config_read_client,cons(nandSim.readClient, nil));
   MemServer#(PhysAddrWidth,64,1) hostDma <- mkMemServerRW(backingStoreMMUConfigIndicationProxy.ifc, hostDmaDebugIndicationProxy.ifc, rcs, cons(nandSim.writeClient, nil), cons(backingStoreMMU,cons(algoMMU,nil)));

   // nandsim mmu0
   MMUConfigIndicationProxy nandsimMMU0ConfigIndicationProxy <- mkMMUConfigIndicationProxy(NandsimMMU0ConfigIndication);
   MMU#(PhysAddrWidth) nandsimMMU0 <- mkMMU(0, False, nandsimMMU0ConfigIndicationProxy.ifc);
   MMUConfigRequestWrapper nandsimMMU0ConfigRequestWrapper <- mkMMUConfigRequestWrapper(NandsimMMU0ConfigRequest, nandsimMMU0.request);
   
   // nandsim memory dma0 server
   DmaDebugIndicationProxy nandsimDma0DebugIndicationProxy <- mkDmaDebugIndicationProxy(NandsimDma0DebugIndication);   
   MemServer#(PhysAddrWidth,64,1) nandsimDma0 <- mkMemServerR(nandsimMMU0ConfigIndicationProxy.ifc, nandsimDma0DebugIndicationProxy.ifc, cons(strstr.haystack_read_clients[0],nil), cons(nandsimMMU0,nil));
   mkConnection(nandsimDma0.masters[0], nandSim.memSlaves[0]);
   
   // nandsim mmu1
   MMUConfigIndicationProxy nandsimMMU1ConfigIndicationProxy <- mkMMUConfigIndicationProxy(NandsimMMU1ConfigIndication);
   MMU#(PhysAddrWidth) nandsimMMU1 <- mkMMU(0, False, nandsimMMU1ConfigIndicationProxy.ifc);
   MMUConfigRequestWrapper nandsimMMU1ConfigRequestWrapper <- mkMMUConfigRequestWrapper(NandsimMMU1ConfigRequest, nandsimMMU1.request);
   
   // nandsim memory dma1 server
   DmaDebugIndicationProxy nandsimDma1DebugIndicationProxy <- mkDmaDebugIndicationProxy(NandsimDma1DebugIndication);   
   MemServer#(PhysAddrWidth,64,1) nandsimDma1 <- mkMemServerR(nandsimMMU1ConfigIndicationProxy.ifc, nandsimDma1DebugIndicationProxy.ifc, cons(strstr.haystack_read_clients[1],nil), cons(nandsimMMU1,nil));
   mkConnection(nandsimDma1.masters[0], nandSim.memSlaves[1]);
   
   Vector#(12,StdPortal) portals;

   portals[0] = nandSimRequestWrapper.portalIfc;
   portals[1] = nandSimIndicationProxy.portalIfc; 

   portals[2] = strstrRequestWrapper.portalIfc;
   portals[3] = strstrIndicationProxy.portalIfc; 
   
   portals[4] = backingStoreMMUConfigRequestWrapper.portalIfc;
   portals[5] = backingStoreMMUConfigIndicationProxy.portalIfc;

   portals[6] = algoMMUConfigRequestWrapper.portalIfc;
   portals[7] = algoMMUConfigIndicationProxy.portalIfc;
   
   portals[8] = nandsimMMU0ConfigRequestWrapper.portalIfc;
   portals[9] = nandsimMMU0ConfigIndicationProxy.portalIfc;

   portals[10] = nandsimMMU0ConfigRequestWrapper.portalIfc;
   portals[11] = nandsimMMU0ConfigIndicationProxy.portalIfc;

   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = hostDma.masters;
   interface leds = default_leds;
      
endmodule : mkConnectalTop
