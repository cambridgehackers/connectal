// bsv libraries
import Vector::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import Portal::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import AxiMasterSlave::*;


// generated by tool
import PortalPerfIndicationProxy::*;
import PortalPerfRequestWrapper::*;

// defined by user
import PortalPerf::*;

typedef enum {PortalPerfIndication, PortalPerfRequest} IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalTop#(addrWidth));

   // instantiate user portals
   PortalPerfIndicationProxy portalperfIndicationProxy <- mkPortalPerfIndicationProxy(PortalPerfIndication);
   PortalPerfRequestWrapper portalperfRequestWrapper <- mkPortalPerfRequestWrapper(PortalPerfRequest);
   
   PortalPerf portalperf <- mkPortalPerf(portalperfIndicationProxy);
   
   Vector#(2,StdPortal) portals;
   portals[0] = portalperfIndicationProxy.portalIfc;
   portals[1] = portalperfRequestWrapper.portalIfc; 

   let interrupt_mux <- mkInterruptMux(portals);
   
   // instantiate system directory
   StdDirectory dir <- mkStdDirectory(portals);
   
   let ctrl_mux <- mkAxiSlaveMuxDbg(dir,portals);
   
   interface interrupt = interrupt_mux;
   interface ctrl = ctrl_mux;
   interface m_axi = null_axi_master;


endmodule : mkPortalTop
