// Copyright (c) 2015 Connectal Project.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
import GetPut::*;
import Connectable::*;

typedef struct {
   Bit#(addrWidth) address;
   Bit#(dataWidth) data;
   Bit#(4)         burstcount;
   Bool            write;
   Bool            sof;
   Bool            eof;
} AvalonMMRequest#(numeric type addrWidth, numeric type dataWidth) deriving (Bits);

typedef struct {
   Bit#(dataWidth) readdata;
} AvalonMMData#(numeric type dataWidth) deriving (Bits);

interface AvalonMMaster#(numeric type addrWidth, numeric type busWidth);
   interface Get#(AvalonMMRequest#(addrWidth, busWidth)) request;
   interface Put#(AvalonMMData#(busWidth)) response;
endinterface

interface AvalonMSlave#(numeric type addrWidth, numeric type busWidth);
   interface Put#(AvalonMMRequest#(addrWidth, busWidth)) request;
   interface Get#(AvalonMMData#(busWidth)) response;
endinterface

instance Connectable#(AvalonMMaster#(addrWidth, dataWidth), AvalonMSlave#(addrWidth, dataWidth));
   module mkConnection#(AvalonMMaster#(addrWidth, dataWidth) m, AvalonMSlave#(addrWidth, dataWidth) s)(Empty);
      mkConnection(m.request, s.request);
      mkConnection(s.response, m.response);
   endmodule
endinstance
