typedef enum {IfcNames_ReadTestIndicationH2S=8, IfcNames_ReadTestRequestS2H} TileNames deriving (Eq,Bits);
