

typedef enum {DmaIndication, DmaConfig, NandSimIndication, NandSimRequest, AlgoIndication, AlgoRequest, NandsimDmaIndication, NandsimDmaConfig} IfcNames deriving (Eq,Bits);

