// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import BlueScope::*;
import PortalMemory::*;
import MemTypes::*;
import DmaUtils::*;
import MemServer::*;
import SGList::*;

// generated by tool
import MaxcommonsubseqRequestWrapper::*;
import DmaDebugRequestWrapper::*;
import SGListConfigRequestWrapper::*;
import MaxcommonsubseqIndicationProxy::*;
import DmaDebugIndicationProxy::*;
import SGListConfigIndicationProxy::*;

// defined by user
import Maxcommonsubseq::*;

typedef enum {MaxcommonsubseqIndication, MaxcommonsubseqRequest, HostmemDmaDebugIndication, HostmemDmaDebugRequest, HostmemSGListConfigRequest, HostmemSGListConfigIndication} IfcNames deriving (Eq,Bits);
typedef 1 DegPar;


module mkPortalTop(StdPortalDmaTop#(PhysAddrWidth));

   DmaReadBuffer#(64,1) setupA_read_chan <- mkDmaReadBuffer();
   DmaReadBuffer#(64,1) setupB_read_chan <- mkDmaReadBuffer();
   DmaWriteBuffer#(64,1) fetch_write_chan <- mkDmaWriteBuffer();
   
   ObjectReadClient#(64) setupA_read_client = setupA_read_chan.dmaClient;
   ObjectReadClient#(64) setupB_read_client = setupB_read_chan.dmaClient;
   ObjectWriteClient#(64) fetch_write_client = fetch_write_chan.dmaClient;
   
   Vector#(2,  ObjectReadClient#(64)) readClients;
   readClients[0] = setupA_read_client;
   readClients[1] = setupB_read_client;

   Vector#(1, ObjectWriteClient#(64)) writeClients;
   writeClients[0] = fetch_write_client;


   SGListConfigIndicationProxy hostmemSGListConfigIndicationProxy <- mkSGListConfigIndicationProxy(HostmemSGListConfigIndication);
   SGListMMU#(PhysAddrWidth) hostmemSGList <- mkSGListMMU(0, True, hostmemSGListConfigIndicationProxy.ifc);
   SGListConfigRequestWrapper hostmemSGListConfigRequestWrapper <- mkSGListConfigRequestWrapper(HostmemSGListConfigRequest, hostmemSGList.request);

   DmaDebugIndicationProxy hostmemDmaDebugIndicationProxy <- mkDmaDebugIndicationProxy(HostmemDmaDebugIndication);
   MemServer#(PhysAddrWidth,64,1) dma <- mkMemServerRW(hostmemDmaDebugIndicationProxy.ifc, readClients, writeClients, hostmemSGList);
   DmaDebugRequestWrapper hostmemDmaDebugRequestWrapper <- mkDmaDebugRequestWrapper(HostmemDmaDebugRequest, dma.request);
   
   MaxcommonsubseqIndicationProxy maxcommonsubseqIndicationProxy <- mkMaxcommonsubseqIndicationProxy(MaxcommonsubseqIndication);
   MaxcommonsubseqRequest maxcommonsubseqRequest <- mkMaxcommonsubseqRequest(maxcommonsubseqIndicationProxy.ifc, setupA_read_chan.dmaServer, setupB_read_chan.dmaServer, fetch_write_chan.dmaServer);
   MaxcommonsubseqRequestWrapper maxcommonsubseqRequestWrapper <- mkMaxcommonsubseqRequestWrapper(MaxcommonsubseqRequest,maxcommonsubseqRequest);

   Vector#(6,StdPortal) portals;
   portals[0] = maxcommonsubseqRequestWrapper.portalIfc;
   portals[1] = maxcommonsubseqIndicationProxy.portalIfc; 
   portals[2] = hostmemDmaDebugRequestWrapper.portalIfc;
   portals[3] = hostmemDmaDebugIndicationProxy.portalIfc; 
   portals[4] = hostmemSGListConfigRequestWrapper.portalIfc;
   portals[5] = hostmemSGListConfigIndicationProxy.portalIfc;

   
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;
endmodule
