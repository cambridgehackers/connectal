// Copyright (c) 2014 Quanta Research Cambridge, Inc.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

// bsv libraries
import Vector::*;
import FIFO::*;
import DefaultValue::*;

// portz libraries
import Portal::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
//import Dma::*;

// generated by tool
import ImageCaptureIndicationProxy::*;
import ImageCaptureRequestWrapper::*;
import ImageonSerdesIndicationProxy::*;
import ImageonSerdesRequestWrapper::*;
import HdmiInternalIndicationProxy::*;
import HdmiInternalRequestWrapper::*;
import ImageonSensorRequestWrapper::*;

// defined by user
import FrequencyCounter::*;
import ImageCapture::*;
import GetPut::*;
import Connectable :: *;
import Clocks :: *;
import XbsvSpi :: *;

import Imageon::*;
import IserdesDatadeser::*;
import HDMI::*;
import XilinxCells::*;
import XbsvXilinxCells::*;
import YUV::*;
//import PS7LIB :: *;
import Imageon :: *;

typedef enum { ImageCapture, ImageonSerdesRequest, HdmiInternalRequest, ImageonSensorRequest,
    ImageCaptureIndication, ImageonSerdesIndication, HdmiInternalIndication} IfcNames deriving (Eq,Bits);

interface ImageCapturePins;
   interface SpiPins spi;
   interface ImageonSensorPins pins;
   interface ImageonSerdesPins serpins;
   interface HDMI hdmi;
   method Bit#(1) i2c_mux_reset_n();
endinterface

module mkPortalTop#(Clock clock200, Clock fmc_imageon_clk1)(PortalTop#(addrWidth,64,ImageCapturePins,0));
   Clock defaultClock <- exposeCurrentClock();
   Reset defaultReset <- exposeCurrentReset();
   IDELAYCTRL idel <- mkIDELAYCTRL(2, clocked_by clock200);
   ClockGenerator7AdvParams clockParams = defaultValue;
   clockParams.bandwidth          = "OPTIMIZED";
   clockParams.compensation       = "ZHOLD";
   clockParams.clkfbout_mult_f    = 8.000;
   clockParams.clkfbout_phase     = 0.0;
   clockParams.clkin1_period      = 6.734007; // 148.5 MHz
   clockParams.clkin2_period      = 6.734007;
   clockParams.clkout0_divide_f   = 8.000;    // 148.5 MHz
   clockParams.clkout0_duty_cycle = 0.5;
   clockParams.clkout0_phase      = 0.0000;
   clockParams.clkout1_divide     = 32;       // 37.125 MHz
   clockParams.clkout1_duty_cycle = 0.5;
   clockParams.clkout1_phase      = 0.0000;
   clockParams.divclk_divide      = 1;
   clockParams.ref_jitter1        = 0.010;
   clockParams.ref_jitter2        = 0.010;

   ClockGenerator7 clockGen <- mkClockGenerator7Adv(clockParams, clocked_by fmc_imageon_clk1);
   Clock hdmi_clock <- mkClockBUFG(clocked_by clockGen.clkout0);    // 148.5   MHz
   Clock imageon_clock <- mkClockBUFG(clocked_by clockGen.clkout1); //  37.125 MHz

   Reset fmc_imageon_reset <- mkAsyncReset(2, defaultReset, fmc_imageon_clk1);
   Reset hdmi_reset <- mkAsyncReset(2, defaultReset, hdmi_clock);
   Reset imageon_reset <- mkAsyncReset(2, defaultReset, imageon_clock);
   SPI#(Bit#(26)) spiController <- mkSPI(1000);
   SyncPulseIfc vsyncPulse <- mkSyncHandshake(hdmi_clock, hdmi_reset, imageon_clock);
   Reg#(Bit#(1)) i2c_mux_reset_n_reg <- mkReg(0);

   // instantiate user portals
   // serdes: serial line protocol for wires from sensor (nothing sensor specific)
   ImageonSerdesIndicationProxy serdesIndicationProxy <- mkImageonSerdesIndicationProxy(ImageonSerdesIndication);
   ISerdes serdes <- mkISerdes(defaultClock, defaultReset, serdesIndicationProxy.ifc,
			clocked_by imageon_clock, reset_by imageon_reset);
   ImageonSerdesRequestWrapper serdesRequestWrapper <- mkImageonSerdesRequestWrapper(ImageonSerdesRequest,serdes.control);

   // hdmi: output to display
   HdmiInternalIndicationProxy hdmiIndicationProxy <- mkHdmiInternalIndicationProxy(HdmiInternalIndication);
   HdmiGenerator hdmiGen <- mkHdmiGenerator(defaultClock, defaultReset,
       vsyncPulse, hdmiIndicationProxy.ifc, clocked_by hdmi_clock, reset_by hdmi_reset);
   HdmiInternalRequestWrapper hdmiRequestWrapper <- mkHdmiInternalRequestWrapper(HdmiInternalRequest,hdmiGen.control);

   // fromSensor: sensor specific processing of serdes input, resulting in pixels
   ImageonSensor fromSensor <- mkImageonSensor(defaultClock, defaultReset, serdes.data, vsyncPulse.pulse(),
       hdmiGen.control, hdmi_clock, hdmi_reset, clocked_by imageon_clock, reset_by imageon_reset);
   ImageonSensorRequestWrapper sensorRequestWrapper <- mkImageonSensorRequestWrapper(ImageonSensorRequest,fromSensor.control);

   ImageCaptureIndicationProxy captureIndicationProxy <- mkImageCaptureIndicationProxy(ImageCaptureIndication);
   FrequencyCounter axiFreqCounter <- mkFrequencyCounter(defaultClock, defaultReset);
   FrequencyCounter hdmiFreqCounter <- mkFrequencyCounter(hdmi_clock, hdmi_reset);
   FrequencyCounter imageonFreqCounter <- mkFrequencyCounter(imageon_clock, imageon_reset);
   FrequencyCounter fmcFreqCounter <- mkFrequencyCounter(fmc_imageon_clk1, fmc_imageon_reset);
   ImageCaptureRequest imageCaptureRequest = (interface ImageCaptureRequest;
      method Action get_debugind();
         captureIndicationProxy.ifc.debugind(fromSensor.control.get_debugind());
      endmethod
      method Action put_spi_request(Bit#(32) v);
         spiController.request.put(truncate(v));
      endmethod
      method Action set_i2c_mux_reset_n(Bit#(1) v);
	 i2c_mux_reset_n_reg <= v;
      endmethod
      method Action measure_axi_clock_period(Bit#(32) cycles_100mhz);
	 axiFreqCounter.start(cycles_100mhz);
      endmethod
      method Action measure_hdmi_clock_period(Bit#(32) cycles_100mhz);
         hdmiFreqCounter.start(cycles_100mhz);
      endmethod
      method Action measure_imageon_clock_period(Bit#(32) cycles_100mhz);
         imageonFreqCounter.start(cycles_100mhz);
      endmethod
      method Action measure_fmc_clock_period(Bit#(32) cycles_100mhz);
         fmcFreqCounter.start(cycles_100mhz);
      endmethod
      endinterface);
   ImageCaptureRequestWrapper captureRequestWrapper <- mkImageCaptureRequestWrapper(ImageCapture, imageCaptureRequest);

   rule spiControllerResponse;
       Bit#(26) v <- spiController.response.get();
       captureIndicationProxy.ifc.spi_response(extend(v));
   endrule

   rule gotAxiClockPeriod;
      let cycles <- axiFreqCounter.elapsedCycles();
      captureIndicationProxy.ifc.axi_clock_period(cycles);
   endrule
   rule gotHdmiClockPeriod;
      let cycles <- hdmiFreqCounter.elapsedCycles();
      captureIndicationProxy.ifc.hdmi_clock_period(cycles);
   endrule
   rule gotImageonClockPeriod;
      let cycles <- imageonFreqCounter.elapsedCycles();
      captureIndicationProxy.ifc.imageon_clock_period(cycles);
   endrule
   rule gotFmcClockPeriod;
      let cycles <- fmcFreqCounter.elapsedCycles();
      captureIndicationProxy.ifc.fmc_clock_period(cycles);
   endrule

   Reg#(Bool) frameStart <- mkReg(False, clocked_by imageon_clock, reset_by imageon_reset);
   Reg#(Bit#(32)) frameCount <- mkReg(0, clocked_by imageon_clock, reset_by imageon_reset);
   SyncFIFOIfc#(Tuple2#(Bit#(2),Bit#(32))) frameStartSynchronizer <- mkSyncFIFO(2, imageon_clock, imageon_reset, defaultClock);

   rule frameStartRule;
       let monitor = fromSensor.monitor();
       Bool fs = unpack(monitor[0]);
       if (fs && !frameStart) begin
	  // start of frame?
	  // need to cross the clock domain
	  frameStartSynchronizer.enq(tuple2(monitor, frameCount));
	  frameCount <= frameCount + 1;
       end
      frameStart <= fs;
   endrule
   rule frameStartIndication;
      let tpl = frameStartSynchronizer.first();
      frameStartSynchronizer.deq();
      let monitor = tpl_1(tpl);
      let count = tpl_2(tpl);
      captureIndicationProxy.ifc.frameStart(monitor, count);
   endrule

   rule xsviConnection;
       // copy data from sensor to hdmi output
       let xsvi <- fromSensor.get_data();
       Bit#(32) pixel = {8'b0, xsvi[9:2], xsvi[9:2], xsvi[9:2]};
       hdmiGen.request.put(pixel);
   endrule
   
   Vector#(7,StdPortal) portals;
   portals[0] = captureRequestWrapper.portalIfc;
   portals[1] = captureIndicationProxy.portalIfc;
   portals[2] = serdesRequestWrapper.portalIfc; 
   portals[3] = serdesIndicationProxy.portalIfc;
   portals[4] = hdmiRequestWrapper.portalIfc; 
   portals[5] = hdmiIndicationProxy.portalIfc; 
   portals[6] = sensorRequestWrapper.portalIfc; 
   
   // instantiate system directory
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = nil;
   //interface leds = captureRequestInternal.leds;

   interface ImageCapturePins pins;
       interface SpiPins spi = spiController.pins;
       interface ImageonSensorPins pins = fromSensor.pins;
       interface ImageonSerdesPins serpins = serdes.pins;
       interface HDMI hdmi = hdmiGen.hdmi;
       method Bit#(1) i2c_mux_reset_n(); return i2c_mux_reset_n_reg; endmethod
   endinterface
endmodule : mkPortalTop
