// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import CtrlMux::*;
import Portal::*;
import Leds::*;
import ConnectalMemory::*;
import MemTypes::*;
import MemServer::*;
import MMU::*;

// generated by tool
import TestRequest::*;
import DmaDebugRequest::*;
import MMUConfigRequest::*;
import TestIndication::*;
import DmaDebugIndication::*;
import MMUConfigIndication::*;

// defined by user
import Test::*;

typedef enum {TestIndication, TestRequest, HostMMUConfigRequest, HostMMUConfigIndication, HostDmaDebugIndication, HostDmaDebugRequest} IfcNames deriving (Eq,Bits);

module mkConnectalTop(StdConnectalDmaTop#(PhysAddrWidth));

   TestIndicationProxy testIndicationProxy <- mkTestIndicationProxy(TestIndication);
   Test test <- mkTestRequest(testIndicationProxy.ifc);
   TestRequestWrapper testRequestWrapper <- mkTestRequestWrapper(TestRequest,test.request);

   MMUConfigIndicationProxy hostMMUConfigIndicationProxy <- mkMMUConfigIndicationProxy(HostMMUConfigIndication);
   MMU#(PhysAddrWidth) hostMMU <- mkMMU(0, True, hostMMUConfigIndicationProxy.ifc);
   MMUConfigRequestWrapper hostMMUConfigRequestWrapper <- mkMMUConfigRequestWrapper(HostMMUConfigRequest, hostMMU.request);

   DmaDebugIndicationProxy hostDmaDebugIndicationProxy <- mkDmaDebugIndicationProxy(HostDmaDebugIndication);
   MemServer#(PhysAddrWidth,64,1) dma <- mkMemServerR(hostMMUConfigIndicationProxy.ifc,
						      hostDmaDebugIndicationProxy.ifc, cons(test.readClient,nil), cons(hostMMU,nil));
   DmaDebugRequestWrapper hostDmaDebugRequestWrapper <- mkDmaDebugRequestWrapper(HostDmaDebugRequest, dma.request);

   Vector#(4,StdPortal) portals;
   portals[0] = testRequestWrapper.portalIfc;
   portals[1] = testIndicationProxy.portalIfc; 
   portals[2] = hostMMUConfigRequestWrapper.portalIfc;
   portals[3] = hostMMUConfigIndicationProxy.portalIfc;
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;
endmodule


