// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import AxiMasterSlave::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import BlueScope::*;
import PortalMemory::*;
import Dma::*;
import DmaUtils::*;
import AxiDma::*;

// generated by tool
import StrstrRequestWrapper::*;
import DmaConfigWrapper::*;
import StrstrIndicationProxy::*;
import DmaIndicationProxy::*;
import DmaDbgIndicationProxy::*;
import DmaDbgConfigWrapper::*;

// defined by user
import Strstr::*;

typedef enum {StrstrIndication, StrstrRequest, DmaIndication, DmaConfig, DmaDbgIndication, DmaDbgConfig} IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalTop#(addrWidth)) 

   provisos(Add#(addrWidth, a__, 52),
	    Add#(b__, addrWidth, 64),
	    Add#(c__, 12, addrWidth),
	    Add#(addrWidth, d__, 44),
	    Add#(e__, c__, 40),
	    Add#(f__, addrWidth, 40));

   DmaIndicationProxy dmaIndicationProxy <- mkDmaIndicationProxy(DmaIndication);
   DmaDbgIndicationProxy dmaDbgIndicationProxy <- mkDmaDbgIndicationProxy(DmaDbgIndication);
   DmaReadBuffer#(64,1) haystack_read_chan <- mkDmaReadBuffer();
   DmaReadBuffer#(64,1) needle_read_chan <- mkDmaReadBuffer();
   DmaReadBuffer#(64,1) mp_next_read_chan <- mkDmaReadBuffer();
   
   Vector#(3, DmaReadClient#(64)) readClients = newVector();
   readClients[0] = haystack_read_chan.dmaClient;
   readClients[1] = needle_read_chan.dmaClient;
   readClients[2] = mp_next_read_chan.dmaClient;

   Vector#(0, DmaWriteClient#(64)) writeClients = newVector();
   Integer numRequests = 8;
   AxiDmaServer#(addrWidth,64) dma <- mkAxiDmaServer(dmaIndicationProxy.ifc, dmaDbgIndicationProxy.ifc, numRequests, readClients, writeClients);
   DmaConfigWrapper dmaConfigWrapper <- mkDmaConfigWrapper(DmaConfig, dma.request);
   DmaDbgConfigWrapper dmaDbgConfigWrapper <- mkDmaDbgConfigWrapper(DmaDbgConfig, dma.dbgRequest);
   
   
   StrstrIndicationProxy strstrIndicationProxy <- mkStrstrIndicationProxy(StrstrIndication);
   StrstrRequest strstrRequest <- mkStrstrRequest(strstrIndicationProxy.ifc, haystack_read_chan.dmaServer, 
						  needle_read_chan.dmaServer, mp_next_read_chan.dmaServer);
   StrstrRequestWrapper strstrRequestWrapper <- mkStrstrRequestWrapper(StrstrRequest,strstrRequest);

   Vector#(6,StdPortal) portals;
   portals[0] = strstrRequestWrapper.portalIfc;
   portals[1] = strstrIndicationProxy.portalIfc; 
   portals[2] = dmaConfigWrapper.portalIfc;
   portals[3] = dmaIndicationProxy.portalIfc; 
   portals[4] = dmaDbgConfigWrapper.portalIfc;
   portals[5] = dmaDbgIndicationProxy.portalIfc;
   
   Directory dir <- mkDirectory(portals);
   Vector#(1,StdPortal) directories;
   directories[0] = dir.portalIfc;
   
   // when constructing ctrl and interrupt muxes, directories must be the first argument
   let ctrl_mux <- mkAxiSlaveMux(directories,portals);
   let interrupt_mux <- mkInterruptMux(portals);
   
   interface interrupt = interrupt_mux;
   interface ctrl = ctrl_mux;
   interface m_axi = dma.m_axi;
   interface leds = default_leds;
endmodule
