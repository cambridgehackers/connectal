// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import AxiMasterSlave::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import BlueScope::*;
import PortalMemory::*;
import PortalRMemory::*;
import AxiDMA::*;

// generated by tool
import StrstrRequestWrapper::*;
import DMARequestWrapper::*;
import StrstrIndicationProxy::*;
import DMAIndicationProxy::*;

// defined by user
import Strstr::*;

typedef enum {StrstrIndication, StrstrRequest, DMAIndication, DMARequest} IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalDmaTop#(addrWidth)) provisos (
    Add#(addrWidth, a__, 52),
    Add#(b__, addrWidth, 64),
    Add#(c__, 12, addrWidth),
    Add#(addrWidth, d__, 44));

   DMAIndicationProxy dmaIndicationProxy <- mkDMAIndicationProxy(DMAIndication);
   DMAReadBuffer#(64,1) haystack_read_chan <- mkDMAReadBuffer();
   DMAReadBuffer#(64,1) needle_read_chan <- mkDMAReadBuffer();
   DMAReadBuffer#(64,1) mp_next_read_chan <- mkDMAReadBuffer();
   
   Vector#(3, DMAReadClient#(64)) readClients = newVector();
   readClients[0] = haystack_read_chan.dmaClient;
   readClients[1] = needle_read_chan.dmaClient;
   readClients[2] = mp_next_read_chan.dmaClient;

   Vector#(0, DMAWriteClient#(64)) writeClients = newVector();
   Integer numRequests = 8;
   AxiDMAServer#(addrWidth,64) dma <- mkAxiDMAServer(dmaIndicationProxy.ifc, numRequests, readClients, writeClients);
   DMARequestWrapper dmaRequestWrapper <- mkDMARequestWrapper(DMARequest,dma.request);

   StrstrIndicationProxy strstrIndicationProxy <- mkStrstrIndicationProxy(StrstrIndication);
   StrstrRequest strstrRequest <- mkStrstrRequest(strstrIndicationProxy.ifc, haystack_read_chan.dmaServer, 
						  needle_read_chan.dmaServer, mp_next_read_chan.dmaServer);
   StrstrRequestWrapper strstrRequestWrapper <- mkStrstrRequestWrapper(StrstrRequest,strstrRequest);

   Vector#(4,StdPortal) portals;
   portals[0] = strstrRequestWrapper.portalIfc;
   portals[1] = strstrIndicationProxy.portalIfc; 
   portals[2] = dmaRequestWrapper.portalIfc;
   portals[3] = dmaIndicationProxy.portalIfc; 
   
   Directory dir <- mkDirectory(portals);
   Vector#(1,StdPortal) directories;
   directories[0] = dir.portalIfc;
   
   // when constructing ctrl and interrupt muxes, directories must be the first argument
   let ctrl_mux <- mkAxiSlaveMux(directories,portals);
   let interrupt_mux <- mkInterruptMux(portals);
   
   interface interrupt = interrupt_mux;
   interface ctrl = ctrl_mux;
   interface m_axi = replicate(dma.m_axi);
   interface leds = ?;
endmodule
