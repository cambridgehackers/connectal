// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import PortalMemory::*;
import Dma::*;
import DmaUtils::*;
import MemServer::*;

// generated by tool
import StrstrRequestWrapper::*;
import DmaConfigWrapper::*;
import StrstrIndicationProxy::*;
import DmaIndicationProxy::*;

// defined by user
import Strstr::*;

typedef enum {StrstrIndication, StrstrRequest, DmaIndication, DmaConfig} IfcNames deriving (Eq,Bits);
typedef 2 DegPar;


module mkPortalTop(StdPortalDmaTop#(addrWidth)) 

   provisos(Add#(addrWidth, a__, 52),
	    Add#(b__, addrWidth, 64),
	    Add#(c__, 12, addrWidth),
	    Add#(addrWidth, d__, 44),
	    Add#(e__, c__, 40),
	    Add#(f__, addrWidth, 40));

   DmaIndicationProxy dmaIndicationProxy <- mkDmaIndicationProxy(DmaIndication);
   Vector#(DegPar,DmaReadBuffer#(64,1)) haystack_read_chans <- replicateM(mkDmaReadBuffer());
   Vector#(DegPar,DmaReadBuffer#(64,1)) needle_read_chans <- replicateM(mkDmaReadBuffer());
   Vector#(DegPar,DmaReadBuffer#(64,1)) mp_next_read_chans <- replicateM(mkDmaReadBuffer());
   
   Vector#(TMul#(3,DegPar), ObjectReadClient#(64)) readClients = newVector();
   for(Integer i = 0; i < valueOf(DegPar); i=i+1) begin
      readClients[(3*i)+0] = haystack_read_chans[i].dmaClient;
      readClients[(3*i)+1] = needle_read_chans[i].dmaClient;
      readClients[(3*i)+2] = mp_next_read_chans[i].dmaClient;
   end

   MemServer#(addrWidth,64,1) dma <- mkMemServerR(dmaIndicationProxy.ifc, readClients);
   DmaConfigWrapper dmaConfigWrapper <- mkDmaConfigWrapper(DmaConfig, dma.request);
   
   function ObjectReadServer#(x) rs(DmaReadBuffer#(x,y) rb);
      return rb.dmaServer;
   endfunction
   
   StrstrIndicationProxy strstrIndicationProxy <- mkStrstrIndicationProxy(StrstrIndication);
   StrstrRequest strstrRequest <- mkStrstrRequest(strstrIndicationProxy.ifc, map(rs,haystack_read_chans), 
						  map(rs,needle_read_chans), map(rs,mp_next_read_chans));
   StrstrRequestWrapper strstrRequestWrapper <- mkStrstrRequestWrapper(StrstrRequest,strstrRequest);

   Vector#(4,StdPortal) portals;
   portals[0] = strstrRequestWrapper.portalIfc;
   portals[1] = strstrIndicationProxy.portalIfc; 
   portals[2] = dmaConfigWrapper.portalIfc;
   portals[3] = dmaIndicationProxy.portalIfc; 
   
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;
endmodule
