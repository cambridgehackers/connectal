// bsv libraries
import Vector::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import Portal::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import AxiMasterSlave::*;
import Dma::*;


// generated by tool
import FibIndicationProxy::*;
import FibRequestWrapper::*;

// defined by user
import Fib::*;

typedef enum {FibIndication, FibRequest} IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalTop#(addrWidth));

   // instantiate user portals
   FibIndicationProxy fibIndicationProxy <- mkFibIndicationProxy(FibIndication);
   FibRequest fibRequest <- mkFibRequest(fibIndicationProxy.ifc);
   FibRequestWrapper fibRequestWrapper <- mkFibRequestWrapper(FibRequest,fibRequestInternal.ifc);
   
   Vector#(2,StdPortal) portals;
   portals[0] = fibIndicationProxy.portalIfc;
   portals[1] = fibRequestWrapper.portalIfc; 
   
   // instantiate system directory
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface master = null_mem_master;
   interface leds = default_leds;

endmodule : mkPortalTop
