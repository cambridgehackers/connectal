/* Copyright (c) 2014 Quanta Research Cambridge, Inc
 *
 * Permission is hereby granted, free of charge, to any person obtaining a
 * copy of this software and associated documentation files (the "Software"),
 * to deal in the Software without restriction, including without limitation
 * the rights to use, copy, modify, merge, publish, distribute, sublicense,
 * and/or sell copies of the Software, and to permit persons to whom the
 * Software is furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included
 * in all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
 * OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
 * FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
 * DEALINGS IN THE SOFTWARE.
 */
import Vector::*;
import FIFO::*;
import GetPut::*;
import Pipe::*;
import Connectable::*;
import CtrlMux::*;
import Portal::*;
import HostInterface::*;
import Leds::*;
import MemPortal::*;
import BlueNoC::*;
import BnocPortal::*;
import BsimLink::*;

// generated by tool
import Simple::*;
import Link::*;

// defined by user
import SimpleIF::*;

typedef enum {SimpleRequest, SimpleIndication, LinkRequest} IfcNames deriving (Eq,Bits);

module mkConnectalTop(StdConnectalTop#(PhysAddrWidth));

   // instantiate user portals
   // the indications from simpleRequest will be connected to the request interface to simpleReuqest2
   SimpleProxyPortal simple1IndicationProxy <- mkSimpleProxyPortal(SimpleIndication);
   Simple simple1 <- mkSimple(simple1IndicationProxy.ifc);
   SimpleWrapper simple1RequestWrapper <- mkSimpleWrapper(SimpleRequest,simple1);

   SimpleProxy simple2IndicationProxy <- mkSimpleProxy(SimpleIndication);
   Simple simple2 <- mkSimple(simple2IndicationProxy.ifc);
   SimpleWrapperPortal simple2RequestWrapper <- mkSimpleWrapperPortal(SimpleRequest, simple2);

   // now connect them via a BlueNoC link
   MsgSource#(4) simpleMsgSource <- mkPortalMsgSource(simple1IndicationProxy.portalIfc);
   MsgSink#(4) simpleMsgSink <- mkPortalMsgSink(simple2RequestWrapper.portalIfc);

   BsimLink link <- mkBsimLink("simplelink");
   (* fire_when_enabled *)
   rule tx;
      simpleMsgSource.dst_rdy(link.tx.notFull());
      if (link.tx.notFull() && simpleMsgSource.src_rdy()) begin
	 let v = simpleMsgSource.beat(); 
	 link.tx.enq(v);
      end
   endrule	    
   (* fire_when_enabled *)
   rule rx;
      simpleMsgSink.src_rdy(link.rx.notEmpty());
      if (link.rx.notEmpty() && simpleMsgSink.dst_rdy()) begin
	 let v <- toGet(link.rx).get();
	 simpleMsgSink.beat(v);
      end
   endrule	    

   Link linkRequest = (interface Link;
		       method Action start(Bool l);
			  link.start(l);
		       endmethod
		       endinterface);
   LinkWrapper linkWrapper <- mkLinkWrapper(LinkRequest, linkRequest);

   Vector#(3,StdPortal) portals;
   portals[0] = simple2IndicationProxy.portalIfc;
   portals[1] = simple1RequestWrapper.portalIfc;
   portals[2] = linkWrapper.portalIfc;
   let ctrl_mux <- mkSlaveMux(portals);

   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = nil;
   interface leds = default_leds;

endmodule : mkConnectalTop
