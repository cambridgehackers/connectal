// bsv libraries
import Vector::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import AxiMasterSlave::*;

// generated by tool
import StructIndicationProxy::*;
import StructRequestWrapper::*;

// defined by user
import Struct::*;

typedef enum {StructIndication, StructRequest} IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalTop#(addrWidth));

   // instantiate user portals
   StructIndicationProxy structIndicationProxy <- mkStructIndicationProxy(StructIndication);
   StructRequest structRequest <- mkStructRequest(structIndicationProxy.ifc);
   StructRequestWrapper structRequestWrapper <- mkStructRequestWrapper(StructRequest,structRequest);
   
   Vector#(2,StdPortal) portals;
   portals[0] = structRequestWrapper.portalIfc; 
   portals[1] = structIndicationProxy.portalIfc;
   let interrupt_mux <- mkInterruptMux(portals);
   
   // instantiate system directory
   StdDirectory dir <- mkStdDirectory(portals);
   Vector#(1,StdPortal) directories;
   directories[0] = dir.portalIfc;
   
   // when constructing the ctrl mux, directories must be the first argument
   let ctrl_mux <- mkAxiSlaveMux(directories,portals);
   
   interface interrupt = interrupt_mux;
   interface ctrl = ctrl_mux;
   interface m_axi = null_axi_master;
   interface leds = default_leds;

endmodule : mkPortalTop


