// Copyright (c) 2013 Quanta Research Cambridge, Inc.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import PortalMemory::*;
import MemTypes::*;
import MemServer::*;
import SGList::*;

// generated by tool
import MemcpyRequestWrapper::*;
import DmaDebugRequestWrapper::*;
import SGListConfigRequestWrapper::*;
import MemcpyIndicationProxy::*;
import DmaDebugIndicationProxy::*;
import SGListConfigIndicationProxy::*;

// defined by user
import Memcpy::*;

typedef enum {MemcpyIndication, 
	      MemcpyRequest, 

	      HostmemDmaDebugIndication, 
	      HostmemDmaDebugRequest, 

	      HostmemSGList0ConfigRequest, 
	      HostmemSGList0ConfigIndication,
	      
	      HostmemSGList1ConfigRequest, 
	      HostmemSGList1ConfigIndication,
	      
	      HostmemSGList2ConfigRequest, 
	      HostmemSGList2ConfigIndication,

	      HostmemSGList3ConfigRequest, 
	      HostmemSGList3ConfigIndication } IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalDmaTop#(PhysAddrWidth));

   MemcpyIndicationProxy memcpyIndicationProxy <- mkMemcpyIndicationProxy(MemcpyIndication);
   Memcpy memcpy <- mkMemcpy(memcpyIndicationProxy.ifc);
   MemcpyRequestWrapper memcpyRequestWrapper <- mkMemcpyRequestWrapper(MemcpyRequest,memcpy.request);


   SGListConfigIndicationProxy hostmemSGList0ConfigIndicationProxy <- mkSGListConfigIndicationProxy(HostmemSGList0ConfigIndication);
   SGListMMU#(PhysAddrWidth) hostmemSGList0 <- mkSGListMMU(0, True, hostmemSGList0ConfigIndicationProxy.ifc);
   SGListConfigRequestWrapper hostmemSGList0ConfigRequestWrapper <- mkSGListConfigRequestWrapper(HostmemSGList0ConfigRequest, hostmemSGList0.request);
   
   SGListConfigIndicationProxy hostmemSGList1ConfigIndicationProxy <- mkSGListConfigIndicationProxy(HostmemSGList1ConfigIndication);
   SGListMMU#(PhysAddrWidth) hostmemSGList1 <- mkSGListMMU(1, True, hostmemSGList1ConfigIndicationProxy.ifc);
   SGListConfigRequestWrapper hostmemSGList1ConfigRequestWrapper <- mkSGListConfigRequestWrapper(HostmemSGList1ConfigRequest, hostmemSGList1.request);
   
   SGListConfigIndicationProxy hostmemSGList2ConfigIndicationProxy <- mkSGListConfigIndicationProxy(HostmemSGList2ConfigIndication);
   SGListMMU#(PhysAddrWidth) hostmemSGList2 <- mkSGListMMU(2, True, hostmemSGList2ConfigIndicationProxy.ifc);
   SGListConfigRequestWrapper hostmemSGList2ConfigRequestWrapper <- mkSGListConfigRequestWrapper(HostmemSGList2ConfigRequest, hostmemSGList2.request);

   SGListConfigIndicationProxy hostmemSGList3ConfigIndicationProxy <- mkSGListConfigIndicationProxy(HostmemSGList3ConfigIndication);
   SGListMMU#(PhysAddrWidth) hostmemSGList3 <- mkSGListMMU(3, True, hostmemSGList3ConfigIndicationProxy.ifc);
   SGListConfigRequestWrapper hostmemSGList3ConfigRequestWrapper <- mkSGListConfigRequestWrapper(HostmemSGList3ConfigRequest, hostmemSGList3.request);
   
   Vector#(1,  ObjectReadClient#(64))   readClients = cons(memcpy.dmaReadClient, nil);
   Vector#(1, ObjectWriteClient#(64))  writeClients = cons(memcpy.dmaWriteClient, nil);

   DmaDebugIndicationProxy hostmemDmaDebugIndicationProxy <- mkDmaDebugIndicationProxy(HostmemDmaDebugIndication);
   let sgls = cons(hostmemSGList0,cons(hostmemSGList1, cons(hostmemSGList2,cons(hostmemSGList3,nil))));  
   MemServer#(PhysAddrWidth,64,1) dma <- mkMemServerRW(hostmemDmaDebugIndicationProxy.ifc, readClients, writeClients, sgls);
   DmaDebugRequestWrapper hostmemDmaDebugRequestWrapper <- mkDmaDebugRequestWrapper(HostmemDmaDebugRequest, dma.request);

   Vector#(12,StdPortal) portals;
   portals[0] = memcpyRequestWrapper.portalIfc;
   portals[1] = memcpyIndicationProxy.portalIfc; 
   portals[2] = hostmemDmaDebugRequestWrapper.portalIfc;
   portals[3] = hostmemDmaDebugIndicationProxy.portalIfc; 
   
   portals[4] = hostmemSGList0ConfigRequestWrapper.portalIfc;
   portals[5] = hostmemSGList0ConfigIndicationProxy.portalIfc;
   
   portals[6] = hostmemSGList1ConfigRequestWrapper.portalIfc;
   portals[7] = hostmemSGList1ConfigIndicationProxy.portalIfc;
   
   portals[8] = hostmemSGList2ConfigRequestWrapper.portalIfc;
   portals[9] = hostmemSGList2ConfigIndicationProxy.portalIfc;

   portals[10] = hostmemSGList3ConfigRequestWrapper.portalIfc;
   portals[11] = hostmemSGList3ConfigIndicationProxy.portalIfc;
   
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;
endmodule


