
// Device Under Test
interface DUT;
    method ActionValue#(Bit#(32)) operate(Bit#(32) a, Bit#(32) b);
endinterface
