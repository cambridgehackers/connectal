// bsv libraries
import Vector::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import Portal::*;
import Directory::*;
import CtrlMux::*;
import Leds::*;
import MemTypes::*;
import HostInterface::*;

// generated by tool
import FpMulIndicationProxy::*;
import FpMulRequestWrapper::*;

// defined by user
import RbmTypes::*;
import FpMacTb::*;

module  mkConnectalTop#(HostType host)(ConnectalTop#(PhysAddrWidth,TMul#(32,N),Empty,NumberOfMasters));

   FpMulIndicationProxy ind <- mkFpMulIndicationProxy(FpMulIndicationPortal);
   FpMulRequest req <- mkFpMulRequest(ind.ifc);
   FpMulRequestWrapper reqW <- mkFpMulRequestWrapper(FpMulRequestPortal,req);

   Vector#(2,StdPortal) portals;
   portals[0] = ind.portalIfc;
   portals[1] = reqW.portalIfc; 
   
   StdDirectory dir <- mkStdDirectory(portals);
   
   // when constructing ctrl and interrupt muxes, directories must be the first argument
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = replicate(?);

endmodule : mkConnectalTop
