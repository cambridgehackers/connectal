// bsv libraries
export Aurora::*;
export mkConnectalTop;

import Vector::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import CtrlMux::*;
import Portal::*;
import Leds::*;
import MemTypes::*;
import MemPortal::*;

// generated by tool
import AuroraIndicationProxy::*;
import AuroraRequestWrapper::*;

// defined by user
import Aurora::*;
typedef enum {AuroraIndication, AuroraRequest} IfcNames deriving (Eq,Bits);

module mkConnectalTop(ConnectalTop#(PhysAddrWidth,64,AuroraPins,0));

   // instantiate user portals
   AuroraIndicationProxy auroraIndicationProxy <- mkAuroraIndicationProxy(AuroraIndication);
   let auroraRequest <- mkAuroraRequest(auroraIndicationProxy.ifc);
   AuroraRequestWrapper auroraRequestWrapper <- mkAuroraRequestWrapper(AuroraRequest,auroraRequest.request);
   
   Vector#(2,StdPortal) portals;
   portals[0] = auroraRequestWrapper.portalIfc;
   portals[1] = auroraIndicationProxy.portalIfc;
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = nil;
   interface leds = default_leds;
   interface pins = auroraRequest.pins;

endmodule : mkConnectalTop
