
import Vector::*;

// libraries
import Directory::*;
import AxiMasterSlave::*;

// generated by tool
import SayWrapper::*;
import SayProxy::*;
import DirectoryRequestWrapper::*;
import DirectoryResponseProxy::*;

// defined by user
import Say::*;

interface Top;
   interface Axi3SlaveStandard ctrl;
   interface Axi3MasterStandard m_axi;      
   interface Vector#(4,ReadOnly#(Bool)) interrupts;
   interface LEDS leds;
endinterface

module mkZynqTop(Top);
   
   Vector#(4, Int) portalMap;
   portalMap[0] = 132;
   portalMap[1] = 56;
   portalMap[2] = 1008;
   portalmap[3] = 7;

   SayProxy sayProxy <- mkSayProxy(7);
   Say say <- mkSay(sayProxy.ifc);
   SayWrapper sayWrapper <- mkSayWrapper(1008,say);
   
   DirectoryResponseProxy dirRespProxy <- mkDirectoryResponseProxy(56)
   DirectoryRequestInternal#(4) dirReqI <- mkDirectoryRequestInternal(dirRespProxy.ifc, portalMap);
   DirectoryRequestWrapper dirReqWrapper <- mkDirectoryRequestWrapper(132,dirReqI.ifc);
   
   Vector#(4,Axi3Slave#(32,32,4,12)) ctrls_v;
   Vector#(4,ReadOnly#(Bool)) interrupts_v;

   ctrls_v[0] = dirReqWrapper.ctrl; // 132
   ctrls_v[1] = dirRespProxy.ctrl;  // 56
   ctrls_v[2] = sayWrapper.ctrl;    // 1008
   ctrls_v[3] = sayProxy.ctrl;      // 7
   let ctrl_mux <- mkAxiSlaveMux(ctrls_v);
   
   interrupts_v[0] = dirWrapper.interrupt;
   interrupts_v[1] = dirRespProxy.interrupt;
   interrupts_v[2] = sayWrapper.interrupt;
   interrupts_v[3] = sayProxy.interrupt;
   
   interface Axi3Master m_axi = ?;
   interface Axi3Slave ctrl = ctrl_mux;
   interface Vector interrupts = interrupt_v;
   interface LEDS leds = ?;
endmodule


import "BDPI" function Action      initPortal(Bit#(32) d);
import "BDPI" function Bool                    writeReq();
import "BDPI" function ActionValue#(Bit#(32)) writeAddr();
import "BDPI" function ActionValue#(Bit#(32)) writeData();
import "BDPI" function Bool                     readReq();
import "BDPI" function ActionValue#(Bit#(32))  readAddr();
import "BDPI" function Action        readData(Bit#(32) d);


module mkBsimTop();
   Top top <- mkZynqTop;
   let wf <- mkPipelineFIFO;
   let init_seq = (action 
		      initPortal(0);
		      initPortal(1);
		      initPortal(2);
		      initPortal(3);
                   endaction);
   let init_fsm <- mkOnce(init_seq);
   rule init_rule;
      init_fsm.start;
   endrule
   rule wrReq (writeReq());
      let wa <- writeAddr;
      let wd <- writeData;
      top.ctrl.write.writeAddr(wa,0,0,0,0,0,0);
      wf.enq(wd);
   endrule
   rule wrData;
      wf.deq;
      top.ctrl.write.writeData(wf.first,0,0,0);
   endrule
   rule rdReq (readReq());
      let ra <- readAddr;
      top.ctrl.read.readAddr(ra,0,0,0,0,0,0);
   endrule
   rule rdResp;
      let rd <- top.ctrl.read.readData;
      readData(rd);
   endrule
endmodule
