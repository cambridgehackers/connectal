// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import BlueScope::*;
import PortalMemory::*;
import MemTypes::*;
import DmaUtils::*;
import MemServer::*;
import MMU::*;

// generated by tool
import MaxcommonsubseqRequestWrapper::*;
import DmaDebugRequestWrapper::*;
import MMUConfigRequestWrapper::*;
import MaxcommonsubseqIndicationProxy::*;
import DmaDebugIndicationProxy::*;
import MMUConfigIndicationProxy::*;

// defined by user
import Maxcommonsubseq::*;

typedef enum {MaxcommonsubseqIndication, MaxcommonsubseqRequest, HostDmaDebugIndication, HostDmaDebugRequest, HostMMUConfigRequest, HostMMUConfigIndication} IfcNames deriving (Eq,Bits);
typedef 1 DegPar;


module mkPortalTop(StdPortalDmaTop#(PhysAddrWidth));

   DmaReadBuffer#(64,1) setupA_read_chan <- mkDmaReadBuffer();
   DmaReadBuffer#(64,1) setupB_read_chan <- mkDmaReadBuffer();
   DmaWriteBuffer#(64,1) fetch_write_chan <- mkDmaWriteBuffer();
   
   ObjectReadClient#(64) setupA_read_client = setupA_read_chan.dmaClient;
   ObjectReadClient#(64) setupB_read_client = setupB_read_chan.dmaClient;
   ObjectWriteClient#(64) fetch_write_client = fetch_write_chan.dmaClient;
   
   Vector#(2,  ObjectReadClient#(64)) readClients;
   readClients[0] = setupA_read_client;
   readClients[1] = setupB_read_client;

   Vector#(1, ObjectWriteClient#(64)) writeClients;
   writeClients[0] = fetch_write_client;


   MMUConfigIndicationProxy hostMMUConfigIndicationProxy <- mkMMUConfigIndicationProxy(HostMMUConfigIndication);
   MMU#(PhysAddrWidth) hostMMU <- mkMMU(0, True, hostMMUConfigIndicationProxy.ifc);
   MMUConfigRequestWrapper hostMMUConfigRequestWrapper <- mkMMUConfigRequestWrapper(HostMMUConfigRequest, hostMMU.request);

   DmaDebugIndicationProxy hostDmaDebugIndicationProxy <- mkDmaDebugIndicationProxy(HostDmaDebugIndication);
   MemServer#(PhysAddrWidth,64,1) dma <- mkMemServerRW(hostDmaDebugIndicationProxy.ifc, readClients, writeClients, cons(hostMMU,nil));
   DmaDebugRequestWrapper hostDmaDebugRequestWrapper <- mkDmaDebugRequestWrapper(HostDmaDebugRequest, dma.request);
   
   MaxcommonsubseqIndicationProxy maxcommonsubseqIndicationProxy <- mkMaxcommonsubseqIndicationProxy(MaxcommonsubseqIndication);
   MaxcommonsubseqRequest maxcommonsubseqRequest <- mkMaxcommonsubseqRequest(maxcommonsubseqIndicationProxy.ifc, setupA_read_chan.dmaServer, setupB_read_chan.dmaServer, fetch_write_chan.dmaServer);
   MaxcommonsubseqRequestWrapper maxcommonsubseqRequestWrapper <- mkMaxcommonsubseqRequestWrapper(MaxcommonsubseqRequest,maxcommonsubseqRequest);

   Vector#(6,StdPortal) portals;
   portals[0] = maxcommonsubseqRequestWrapper.portalIfc;
   portals[1] = maxcommonsubseqIndicationProxy.portalIfc; 
   portals[2] = hostDmaDebugRequestWrapper.portalIfc;
   portals[3] = hostDmaDebugIndicationProxy.portalIfc; 
   portals[4] = hostMMUConfigRequestWrapper.portalIfc;
   portals[5] = hostMMUConfigIndicationProxy.portalIfc;

   
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;
endmodule
