
module B2C(C, R, BC, BR);

output C;
output R;
input BC;
input BR;

assign C = BC;
assign R = BR;
endmodule
