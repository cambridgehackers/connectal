typedef enum {ReadTestIndicationH2S=8, ReadTestRequestS2H} TileNames deriving (Eq,Bits);
