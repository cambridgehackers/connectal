// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import AxiMasterSlave::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import PortalMemory::*;
import Dma::*;
import DmaUtils::*;
import PhysicalDma::*;

// generated by tool
import Memread2RequestWrapper::*;
import DmaConfigWrapper::*;
import Memread2IndicationProxy::*;
import DmaIndicationProxy::*;

// defined by user
import Memread2::*;

typedef enum {Memread2Indication, Memread2Request, DmaIndication, DmaConfig} IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalTop#(addrWidth)) provisos (
    Add#(addrWidth, a__, 52),
    Add#(b__, addrWidth, 64),
    Add#(c__, 12, addrWidth),
    Add#(addrWidth, d__, 44),
    Add#(e__, addrWidth, 40),
    Add#(f__, c__, 40));

   DmaIndicationProxy dmaIndicationProxy <- mkDmaIndicationProxy(DmaIndication);

   Memread2IndicationProxy memreadIndicationProxy <- mkMemread2IndicationProxy(Memread2Indication);
   Memread2 memread <- mkMemread2(memreadIndicationProxy.ifc);
   Memread2RequestWrapper memreadRequestWrapper <- mkMemread2RequestWrapper(Memread2Request,memread.request);

   Vector#(2, DmaReadClient#(64)) clients;
   Bool buffered = True;
   if (buffered) begin
      Vector#(2, DmaReadBuffer#(64, 16)) readBuffers <- replicateM(mkDmaReadBuffer);
      mkConnection(memread.dmaClient, readBuffers[0].dmaServer);
      mkConnection(memread.dmaClient2, readBuffers[1].dmaServer);
      clients = cons(readBuffers[0].dmaClient, cons(readBuffers[1].dmaClient, nil));
   end
   else begin
      clients = cons(memread.dmaClient, cons(memread.dmaClient2, nil));
   end

   PhysicalDmaServer#(addrWidth,64) dma <- mkPhysicalDmaServer(dmaIndicationProxy.ifc, clients, nil);

   DmaConfigWrapper dmaRequestWrapper <- mkDmaConfigWrapper(DmaConfig,dma.request);

   Vector#(4,StdPortal) portals;
   portals[0] = memreadRequestWrapper.portalIfc;
   portals[1] = memreadIndicationProxy.portalIfc; 
   portals[2] = dmaRequestWrapper.portalIfc;
   portals[3] = dmaIndicationProxy.portalIfc; 
   
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkAxiSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface ctrl = ctrl_mux;
   interface read_client = dma.read_client;
   interface write_client = dma.write_client;
   interface leds = ?;
endmodule : mkPortalTop
