// Copyright (c) 2016 Accelerated Tech, Inc.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

import Strstr::*;
import Vector::*;
import BuildVector::*;

import ConnectalMemTypes::*;

interface StrstrExample;
   interface StrstrRequest request;
   interface Vector#(2, MemReadClient#(64)) readClients;
endinterface

module mkStrstrExample#(StrstrIndication ind)(StrstrExample);
   Strstr#(64,64) strstr <- mkStrstr(ind);
   interface request = strstr.request;
   interface readClients = append(strstr.config_read_client, strstr.haystack_read_client);
endmodule
