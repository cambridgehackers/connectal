// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import CtrlMux::*;
import Portal::*;
import Leds::*;
import ConnectalMemory::*;
import MemTypes::*;
import MemServer::*;
import MMU::*;

// generated by tool
import MemlatencyRequest::*;
import MemServerRequest::*;
import MMURequest::*;
import MemlatencyIndication::*;
import MemServerIndication::*;
import MMUIndication::*;

// defined by user
import Memlatency::*;

typedef enum {MemlatencyIndication, MemlatencyRequest, HostMemServerIndication, HostMemServerRequest, HostMMURequest, HostMMUIndication} IfcNames deriving (Eq,Bits);

module mkConnectalTop(StdConnectalDmaTop#(PhysAddrWidth));

   MemlatencyIndicationProxy memlatencyIndicationProxy <- mkMemlatencyIndicationProxy(MemlatencyIndication);
   Memlatency memlatency <- mkMemlatency(memlatencyIndicationProxy.ifc);
   MemlatencyRequestWrapper memlatencyRequestWrapper <- mkMemlatencyRequestWrapper(MemlatencyRequest,memlatency.request);
   
   Vector#(1,  MemReadClient#(64))   readClients = cons(memlatency.dmaReadClient, nil);
   Vector#(1, MemWriteClient#(64)) writeClients = cons(memlatency.dmaWriteClient, nil);
   MMUIndicationProxy hostMMUIndicationProxy <- mkMMUIndicationProxy(HostMMUIndication);
   MMU#(PhysAddrWidth) hostMMU <- mkMMU(0, True, hostMMUIndicationProxy.ifc);
   MMURequestWrapper hostMMURequestWrapper <- mkMMURequestWrapper(HostMMURequest, hostMMU.request);

   MemServerIndicationProxy hostMemServerIndicationProxy <- mkMemServerIndicationProxy(HostMemServerIndication);
   MemServer#(PhysAddrWidth,64,1) dma <- mkMemServerRW(hostMemServerIndicationProxy.ifc, readClients, writeClients, cons(hostMMU,nil));
   MemServerRequestWrapper hostMemServerRequestWrapper <- mkMemServerRequestWrapper(HostMemServerRequest, dma.request);
   
   Vector#(6,StdPortal) portals;
   portals[0] = memlatencyRequestWrapper.portalIfc;
   portals[1] = memlatencyIndicationProxy.portalIfc; 
   portals[2] = hostMemServerRequestWrapper.portalIfc;
   portals[3] = hostMemServerIndicationProxy.portalIfc; 
   portals[4] = hostMMURequestWrapper.portalIfc;
   portals[5] = hostMMUIndicationProxy.portalIfc;
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface Empty pins; endinterface
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;
endmodule


