// Copyright (c) 2015 The Connectal Project

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
//import Clocks::*;

interface Clai;
    method Action      deq(Bit#(1) ff);
    //method Bit#(1)     RDY_deq();
    method Action      enq(Bit#(32) v);
    method Bit#(32)    first();
    method Bit#(1)     first__guard();
    method Bit#(1)     notempty();
    method Bit#(1)     notfull();
endinterface

import "BVI" l_class_OC_Fifo1 =
module mkClai(Clai);
    default_clock clk(CLK);
    default_reset rst(RST);
    method deq(deq) enable(EN_deq) ready(RDY_deq);
    method enq(enq_v) enable(enq_ENA);// ready(enq__guard);
    method first first();
    method first__guard first__guard();
    method notEmpty notempty();
    method notFull notfull();
    schedule(first, first__guard, notempty, notfull, deq, enq)
          CF(first, first__guard, notempty, notfull, deq, enq);
endmodule

