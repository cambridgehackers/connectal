
module B2C(B, C);

input B;
output C;

assign C = B;
endmodule
