/* Copyright (c) 2014 Quanta Research Cambridge, Inc
 *
 * Permission is hereby granted, free of charge, to any person obtaining a
 * copy of this software and associated documentation files (the "Software"),
 * to deal in the Software without restriction, including without limitation
 * the rights to use, copy, modify, merge, publish, distribute, sublicense,
 * and/or sell copies of the Software, and to permit persons to whom the
 * Software is furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included
 * in all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
 * OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
 * FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
 * DEALINGS IN THE SOFTWARE.
 */
import Vector::*;
import FIFO::*;
import Connectable::*;
import CtrlMux::*;
import Portal::*;
import HostInterface::*;
import Leds::*;
import MMU::*;
import MemServer::*;
import MemPortal::*;
import SharedMemoryPortal::*;

// generated by tool
import Simple::*;
import MMURequest::*;
import MMUIndication::*;
import SharedMemoryPortalConfig::*;
import MemServerIndication::*;

// defined by user
import SimpleIF::*;

typedef enum {SimpleIndication, SimpleRequest,
	      MMURequest, MMUIndication, MemServerIndication, ReqConfigWrapper, IndConfigWrapper} IfcNames deriving (Eq,Bits);

module mkConnectalTop(StdConnectalDmaTop#(PhysAddrWidth));
   // instantiate DUT
   SimpleProxyPortal indProxy <- mkSimpleProxyPortal(SimpleIndication);
   Simple reqDUT <- mkSimple(indProxy.ifc);
   SimpleWrapperPortal reqWrap <- mkSimpleWrapperPortal(SimpleRequest,reqDUT);
   
   // Use shared memory for DUT requests
   SharedMemoryPortal#(64) reqPortal <- mkSharedMemoryPortal(reqWrap.portalIfc);
   SharedMemoryPortalConfigWrapper reqConfig <-
       mkSharedMemoryPortalConfigWrapper(ReqConfigWrapper, reqPortal.cfg);

   // Use shared memory for DUT indications
   SharedMemoryPortal#(64) indPortal <- mkSharedMemoryPortal(indProxy.portalIfc);
   SharedMemoryPortalConfigWrapper indConfig <-
       mkSharedMemoryPortalConfigWrapper(IndConfigWrapper, indPortal.cfg);

   // MMU used for shared memory buffer mapping
   MMUIndicationProxy indMMU <- mkMMUIndicationProxy(MMUIndication);
   MMU#(PhysAddrWidth) mmu <- mkMMU(0, True, indMMU.ifc);
   MMURequestWrapper reqMMU <- mkMMURequestWrapper(MMURequest, mmu.request);

   let readClients = cons(reqPortal.readClient,
                     cons(indPortal.readClient, nil));
   let writeClients = cons(reqPortal.writeClient,
                      cons(indPortal.writeClient, nil));
   // MemServer used for shared memory buffer access
   MemServerIndicationProxy indMem <- mkMemServerIndicationProxy(MemServerIndication);
   MemServer#(PhysAddrWidth,64,1) dma <- mkMemServerRW(indMem.ifc, readClients, writeClients, cons(mmu,nil));

   Vector#(5,StdPortal) portals;
   portals[0] = reqMMU.portalIfc;
   portals[1] = indMMU.portalIfc;
   portals[2] = reqConfig.portalIfc;
   portals[3] = indConfig.portalIfc;
   portals[4] = indMem.portalIfc;
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;
endmodule : mkConnectalTop
