
/*
   /home/jamey/connectal/generated/scripts/importbvi.py
   -o
   VaddBvi.bsv
   -P
   VaddBvi
   -I
   VaddBvi
   -c
   ap_clk
   -r
   ap_rst
   verilog/vectoradd.v
   -n
   in0
   -n
   in1
   -n
   out
   -n
   ap
*/

import Clocks::*;
import DefaultValue::*;
import XilinxCells::*;
import GetPut::*;
import AxiBits::*;

(* always_ready, always_enabled *)
interface VaddBvi;
    method Bit#(1)     ap_done();
    method Bit#(1)     ap_idle();
    method Bit#(1)     ap_ready();
    method Action      ap_start(Bit#(1) v);
    method Action      in0(Bit#(32) v);
    method Bit#(1)     in0_ap_ack();
    method Action      in0_ap_vld(Bit#(1) v);
    method Action      in1(Bit#(32) v);
    method Bit#(1)     in1_ap_ack();
    method Action      in1_ap_vld(Bit#(1) v);
    method Bit#(32)     out_r();
    method Action      out_r_ap_ack(Bit#(1) v);
    method Bit#(1)     out_r_ap_vld();
endinterface
import "BVI" vectoradd =
module mkVaddBvi(VaddBvi);
   Clock ap_clk <- exposeCurrentClock;
   Reset reset <- exposeCurrentReset;
   Reset ap_rst <- mkResetInverter(reset);
    default_clock ap_clk(ap_clk) = ap_clk;
    default_reset ap_rst(ap_rst) = ap_rst;
    method ap_done ap_done();
    method ap_idle ap_idle();
    method ap_ready ap_ready();
    method ap_start(ap_start) enable((*inhigh*) EN_ap_start);
    method in0(in0) enable((*inhigh*) EN_in0);
    method in0_ap_ack in0_ap_ack();
    method in0_ap_vld(in0_ap_vld) enable((*inhigh*) EN_in0_ap_vld);
    method in1(in1) enable((*inhigh*) EN_in1);
    method in1_ap_ack in1_ap_ack();
    method in1_ap_vld(in1_ap_vld) enable((*inhigh*) EN_in1_ap_vld);
    method out_r out_r();
    method out_r_ap_ack(out_r_ap_ack) enable((*inhigh*) EN_out_r_ap_ack);
    method out_r_ap_vld out_r_ap_vld();
    schedule (ap_done, ap_idle, ap_ready, ap_start, in0, in0_ap_ack, in0_ap_vld, in1, in1_ap_ack, in1_ap_vld, out_r, out_r_ap_ack, out_r_ap_vld) CF (ap_done, ap_idle, ap_ready, ap_start, in0, in0_ap_ack, in0_ap_vld, in1, in1_ap_ack, in1_ap_vld, out_r, out_r_ap_ack, out_r_ap_vld);
endmodule
