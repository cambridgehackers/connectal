// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;


// portz libraries
import AxiMasterSlave::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import PortalMemory::*;
import BlueScope::*;
import AxiRDMA::*;
import BsimRDMA::*;
import PortalMemory::*;
import PortalRMemory::*;
import Directory::*;

// generated by tool
import DirectoryRequestWrapper::*;
import DirectoryResponseProxy::*;
import MemcpyRequestWrapper::*;
import BlueScopeRequestWrapper::*;
import DMARequestWrapper::*;
import MemcpyIndicationProxy::*;
import BlueScopeIndicationProxy::*;
import DMAIndicationProxy::*;

// defined by user
import Memcpy::*;

interface Top;
   interface StdAxi3Slave     ctrl;
   interface StdAxi3Master    m_axi;
   interface ReadOnly#(Bool)  interrupt;
   interface LEDS             leds;
endinterface

module mkZynqTop(Top);

   DMAIndicationProxy dmaIndicationProxy <- mkDMAIndicationProxy(9);
`ifdef BSIM
   BsimDMA#(Bit#(64))  dma <- mkBsimDMA(dmaIndicationProxy.ifc);
`else
   AxiDMA#(Bit#(64))   dma <- mkAxiDMA(dmaIndicationProxy.ifc);
`endif
   DMARequestWrapper dmaRequestWrapper <- mkDMARequestWrapper(1005,dma.request);

   // dma read channel 0 is reserved for memcpy read path
   ReadChan#(Bit#(64)) dma_stream_read_chan = dma.read.readChannels[0];
   // dma write channel 0 is reserved for memcpy write path
   WriteChan#(Bit#(64)) dma_stream_write_chan = dma.write.writeChannels[0];
   // dma read channel 1 is reserved for debug read path
   ReadChan#(Bit#(64)) dma_word_read_chan = dma.read.readChannels[1];
   // dma write channel 1 is reserved for Bluescope output
   WriteChan#(Bit#(64)) dma_debug_write_chan = dma.write.writeChannels[1];

   BlueScopeIndicationProxy blueScopeIndicationProxy <- mkBlueScopeIndicationProxy(8);
   BlueScopeInternal bsi <- mkBlueScopeInternal(32, dma_debug_write_chan, blueScopeIndicationProxy.ifc);
   BlueScopeRequestWrapper blueScopeRequestWrapper <- mkBlueScopeRequestWrapper(1003,bsi.requestIfc);

   MemcpyIndicationProxy memcpyIndicationProxy <- mkMemcpyIndicationProxy(7);
   MemcpyRequest memcpyRequest <- mkMemcpyRequest(memcpyIndicationProxy.ifc, dma_stream_read_chan, dma_stream_write_chan,dma_word_read_chan,bsi);
   MemcpyRequestWrapper memcpyRequestWrapper <- mkMemcpyRequestWrapper(1008,memcpyRequest);

   Vector#(6,StdPortal) portals;
   portals[0] = memcpyRequestWrapper.portalIfc;
   portals[1] = memcpyIndicationProxy.portalIfc; 
   portals[2] = blueScopeRequestWrapper.portalIfc;
   portals[3] = blueScopeIndicationProxy.portalIfc; 
   portals[4] = dmaRequestWrapper.portalIfc;
   portals[5] = dmaIndicationProxy.portalIfc; 
   
   // instantiate system directories
   DirectoryResponseProxy dirRespProxy <- mkDirectoryResponseProxy(56);
   DirectoryRequest dirReq <- mkDirectoryRequest(portals, dirRespProxy.ifc);
   DirectoryRequestWrapper dirReqWrapper <- mkDirectoryRequestWrapper(132,dirReq);

   Vector#(2,StdPortal) directories;
   directories[0] = dirReqWrapper.portalIfc;
   directories[1] = dirRespProxy.portalIfc;
   
   // when constructing ctrl and interrupt muxes, directories must be the first argument
   let ctrl_mux <- mkAxiSlaveMux(directories,portals);
   let interrupt_mux <- mkInterruptMux(directories,portals);
   let axi_master <- mkAxi3Master(dma.m_axi);
   
   interface Vector interrupt = interrupt_mux;
   interface StdAxi3Slave ctrl = ctrl_mux;
`ifndef BSIM
   interface StdAxi3Master m_axi = axi_master;
`endif
endmodule
