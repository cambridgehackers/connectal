
// Copyright (c) 2013 Nokia, Inc.
// Copyright (c) 2013 Quanta Research Cambridge, Inc.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

import FIFO::*;
import SPI::*;

import Zynq::*;
import Imageon::*;
import HDMI::*;

interface ImageCaptureIndications;
endinterface

interface ImageCapture;
    interface ImageonVita imageon;
//    interface HDMI hdmi;
endinterface

module mkImageCapture#(//Clock hdmi_clock, 
       ImageCaptureIndications indications)(ImageCapture);
    interface ImageonVita imageon;
	method Bit#(1) reset_n();
	    return 1;
	endmethod
	method Bit#(3) trigger();
	    return 0;
	endmethod
	method Action monitor(Bit#(2) m);
	endmethod
	method Action data(Bit#(1) sync, Bit#(8) d);
	endmethod
	interface SPI_Pins spiPins;
	endinterface
    endinterface
    // interface HDMI hdmi;
    // 	method Bit#(1) hdmi_vsync;
    // 	    return 0;
    // 	endmethod
    // 	method Bit#(1) hdmi_hsync;
    // 	    return 0;
    // 	endmethod
    // 	method Bit#(1) hdmi_de;
    // 	    return 0;
    // 	endmethod
    // 	method Bit#(16) hdmi_data;
    // 	    return 16'hab;
    // 	endmethod
    // endinterface
endmodule
