// bsv libraries
import Vector::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import Portal::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import AxiMasterSlave::*;


// generated by tool
import BscanIndicationProxy::*;
import BscanRequestWrapper::*;

// defined by user
import BscanRequest::*;

typedef enum {BscanIndication, BscanRequest} IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalTop#(addrWidth));

   // instantiate user portals
   BscanIndicationProxy bscanIndicationProxy <- mkBscanIndicationProxy(BscanIndication);
   BscanRequest bscanRequest <- mkBscanRequest(bscanIndicationProxy.ifc);
   BscanRequestWrapper bscanRequestWrapper <- mkBscanRequestWrapper(BscanRequest,bscanRequest);
   
   Vector#(2,StdPortal) portals;
   portals[0] = bscanIndicationProxy.portalIfc;
   portals[1] = bscanRequestWrapper.portalIfc; 
   let interrupt_mux <- mkInterruptMux(portals);
   
   // instantiate system directory
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkAxiSlaveMux(dir,portals);
   
   interface interrupt = interrupt_mux;
   interface ctrl = ctrl_mux;
   interface m_axi = null_axi_master;

endmodule : mkPortalTop
