// bsv libraries
import Vector::*;
import FIFO::*;
import Connectable::*;
import DefaultValue::*;

// portz libraries
import Portal::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import Dma::*;

// generated by tool
import ImageCaptureIndicationProxy::*;
import ImageCaptureRequestWrapper::*;
import ImageonSerdesIndicationProxy::*;
import HdmiInternalIndicationProxy::*;
//import ImageCaptureRequestInternal::*;
import ImageonSerdesRequestWrapper::*;
import HdmiInternalRequestWrapper::*;
import ImageonSensorRequestWrapper::*;
import ImageCaptureRequestWrapper::*;

// defined by user
import FrequencyCounter::*;
import ImageCapture::*;
import GetPut::*;
import Connectable :: *;
import PCIE :: *; // ConnectableWithClocks
import Clocks :: *;
import XbsvSpi :: *;

import GetPutWithClocks :: *;
import Imageon::*;
import IserdesDatadeser::*;
import HDMI::*;
import SensorToVideo::*;
import XilinxCells::*;
import XbsvXilinxCells::*;
import YUV::*;
import PS7LIB :: *;
import Imageon :: *;

typedef enum { ImageCapture, ImageonSerdesRequest, HdmiInternalRequest, ImageonSensorRequest,
    ImageCaptureIndication, ImageonSerdesIndication, HdmiInternalIndication} IfcNames deriving (Eq,Bits);

interface ImageCapturePins;
   interface SpiPins spi;
   interface ImageonSensorPins pins;
   //interface ImageonTopPins toppins;
   interface ImageonSerdesPins serpins;
   method Bit#(1) i2c_mux_reset_n();
endinterface

module mkPortalTop#(Clock clock200, Clock fmc_imageon_clk1)(PortalTop#(addrWidth,64,ImageCapturePins));
   Clock defaultClock <- exposeCurrentClock();
   Reset defaultReset <- exposeCurrentReset();

   // instantiate user portals
   ImageCaptureIndicationProxy captureIndicationProxy <- mkImageCaptureIndicationProxy(ImageCaptureIndication);
   ImageonSerdesIndicationProxy serdesIndicationProxy <- mkImageonSerdesIndicationProxy(ImageonSerdesIndication);
   HdmiInternalIndicationProxy hdmiIndicationProxy <- mkHdmiInternalIndicationProxy(HdmiInternalIndication);

   //ImageCaptureRequest captureRequestInternal <- mkImageCaptureRequest(captureIndicationProxy.ifc);

//////
   Clock clock200_buf <- mkClockBUFG(clocked_by clock200);
   IDELAYCTRL idel <- mkIDELAYCTRL(2, clocked_by clock200_buf);

   ClockGenerator7AdvParams clockParams = defaultValue;
   clockParams.bandwidth          = "OPTIMIZED";
   clockParams.compensation       = "ZHOLD";
   clockParams.clkfbout_mult_f    = 8.000;
   clockParams.clkfbout_phase     = 0.0;
   clockParams.clkin1_period      = 6.734007; // 148.5 MHz
   clockParams.clkin2_period      = 6.734007;
   clockParams.clkout0_divide_f   = 8.000;    // 148.5 MHz
   clockParams.clkout0_duty_cycle = 0.5;
   clockParams.clkout0_phase      = 0.0000;
   clockParams.clkout1_divide     = 32;       // 37.125 MHz
   clockParams.clkout1_duty_cycle = 0.5;
   clockParams.clkout1_phase      = 0.0000;
   clockParams.divclk_divide      = 1;
   clockParams.ref_jitter1        = 0.010;
   clockParams.ref_jitter2        = 0.010;

   ClockGenerator7 clockGen <- mkClockGenerator7Adv(clockParams, clocked_by fmc_imageon_clk1);
   Clock hdmi_clock = clockGen.clkout0;    // 148.5   MHz
   Clock imageon_clock = clockGen.clkout1; //  37.125 MHz

    Reset fmc_imageon_reset <- mkAsyncReset(2, defaultReset, fmc_imageon_clk1);
    Reset hdmi_reset <- mkAsyncReset(2, defaultReset, hdmi_clock);
    Reset imageon_reset <- mkAsyncReset(2, defaultReset, imageon_clock);
    SyncPulseIfc vsyncPulse <- mkSyncHandshake(hdmi_clock, hdmi_reset, imageon_clock);

    ISerdes serdes <- mkISerdes(defaultClock, defaultReset, serdesIndicationProxy.ifc,
				clocked_by imageon_clock, reset_by imageon_reset);
    SPI#(Bit#(26)) spiController <- mkSPI(1000);
    SensorToVideo converter <- mkSensorToVideo(clocked_by hdmi_clock, reset_by hdmi_reset);
    HdmiGenerator hdmiGen <- mkHdmiGenerator(defaultClock, defaultReset,
        vsyncPulse, hdmiIndicationProxy.ifc, clocked_by hdmi_clock, reset_by hdmi_reset);
    ImageonSensor fromSensor <- mkImageonSensor(defaultClock, defaultReset, serdes.data, vsyncPulse.pulse(),
        hdmiGen.control, hdmi_clock, hdmi_reset, clocked_by imageon_clock, reset_by imageon_reset);

    rule spiControllerResponse;
        Bit#(26) v <- spiController.response.get();
       captureIndicationProxy.ifc.spi_response(extend(v));
    endrule

   Reg#(Bit#(1)) i2c_mux_reset_n_reg <- mkReg(0);
   FrequencyCounter axiFreqCounter <- mkFrequencyCounter(defaultClock, defaultReset);
   FrequencyCounter hdmiFreqCounter <- mkFrequencyCounter(hdmi_clock, hdmi_reset);
   FrequencyCounter imageonFreqCounter <- mkFrequencyCounter(imageon_clock, imageon_reset);
   FrequencyCounter fmcFreqCounter <- mkFrequencyCounter(fmc_imageon_clk1, fmc_imageon_reset);

   rule gotAxiClockPeriod;
      let cycles <- axiFreqCounter.elapsedCycles();
      captureIndicationProxy.ifc.axi_clock_period(cycles);
   endrule
   rule gotHdmiClockPeriod;
      let cycles <- hdmiFreqCounter.elapsedCycles();
      captureIndicationProxy.ifc.hdmi_clock_period(cycles);
   endrule
   rule gotImageonClockPeriod;
      let cycles <- imageonFreqCounter.elapsedCycles();
      captureIndicationProxy.ifc.imageon_clock_period(cycles);
   endrule
   rule gotFmcClockPeriod;
      let cycles <- fmcFreqCounter.elapsedCycles();
      captureIndicationProxy.ifc.fmc_clock_period(cycles);
   endrule

   ImageCaptureRequest imageCaptureRequest = (interface ImageCaptureRequest;
      method Action get_debugind();
         captureIndicationProxy.ifc.debugind(fromSensor.control.get_debugind());
      endmethod
      method Action put_spi_request(Bit#(32) v);
         spiController.request.put(truncate(v));
      endmethod
      method Action set_i2c_mux_reset_n(Bit#(1) v);
	 i2c_mux_reset_n_reg <= v;
      endmethod
      method Action measure_axi_clock_period(Bit#(32) cycles_100mhz);
	 axiFreqCounter.start(cycles_100mhz);
      endmethod
      method Action measure_hdmi_clock_period(Bit#(32) cycles_100mhz);
         hdmiFreqCounter.start(cycles_100mhz);
      endmethod
      method Action measure_imageon_clock_period(Bit#(32) cycles_100mhz);
         imageonFreqCounter.start(cycles_100mhz);
      endmethod
      method Action measure_fmc_clock_period(Bit#(32) cycles_100mhz);
         fmcFreqCounter.start(cycles_100mhz);
      endmethod
      endinterface);

    ImageCaptureRequestWrapper captureRequestWrapper <- mkImageCaptureRequestWrapper(ImageCapture, imageCaptureRequest);
    ImageonSerdesRequestWrapper serdesRequestWrapper <- mkImageonSerdesRequestWrapper(ImageonSerdesRequest,serdes.control);
    HdmiInternalRequestWrapper hdmiRequestWrapper <- mkHdmiInternalRequestWrapper(HdmiInternalRequest,hdmiGen.control);
    ImageonSensorRequestWrapper sensorRequestWrapper <- mkImageonSensorRequestWrapper(ImageonSensorRequest,fromSensor.control);

    rule xsviConnection;
        let xsvi <- fromSensor.get_data();
        //bsi.dataIn(extend(pack(xsvi)), extend(pack(xsvi)));
        //converter.in.put(xsvi);
        //let xvideo <- converter.out.get();
        //hdmiGen.rgb(xvideo);
        Bit#(64) pixel = {40'b0, xsvi[9:2], xsvi[9:2], xsvi[9:2]};
        hdmiGen.request.put(pixel);
    endrule
   
   Vector#(7,StdPortal) portals;
   portals[0] = captureRequestWrapper.portalIfc;
   portals[1] = captureIndicationProxy.portalIfc;
   portals[2] = serdesRequestWrapper.portalIfc; 
   portals[3] = serdesIndicationProxy.portalIfc;
   portals[4] = hdmiRequestWrapper.portalIfc; 
   portals[5] = hdmiIndicationProxy.portalIfc; 
   portals[6] = sensorRequestWrapper.portalIfc; 
   
   // instantiate system directory
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface master = null_mem_master;
   //interface leds = captureRequestInternal.leds;

   interface ImageCapturePins pins;
       interface SpiPins spi = spiController.pins;
       interface ImageonSensorPins pins = fromSensor.pins;
       interface ImageonSerdesPins serpins = serdes.pins;
       method Bit#(1) i2c_mux_reset_n(); return i2c_mux_reset_n_reg; endmethod
   endinterface

endmodule : mkPortalTop
