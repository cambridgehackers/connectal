// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import AxiClientServer::*;
import AxiMasterSlave::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import BlueScope::*;
import PortalMemory::*;
import PortalRMemory::*;
`ifdef BSIM
import BsimRDMA::*;
`else
import AxiRDMA::*;
`endif

// generated by tool
import StrstrRequestWrapper::*;
import DMARequestWrapper::*;
import StrstrIndicationProxy::*;
import DMAIndicationProxy::*;

// defined by user
import Strstr::*;

typedef enum {StrstrIndication, StrstrRequest, DMAIndication, DMARequest} IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalDmaTop);

   DMAIndicationProxy dmaIndicationProxy <- mkDMAIndicationProxy(DMAIndication);
   DMAReadBuffer#(64,8) haystack_read_chan <- mkDMAReadBuffer();
   DMAReadBuffer#(64,8) needle_read_chan <- mkDMAReadBuffer();
   DMAReadBuffer#(64,8) mp_next_read_chan <- mkDMAReadBuffer();
   
   Vector#(3, DMAReadClient#(64)) readClients = newVector();
   readClients[0] = haystack_read_chan.dmaClient;
   readClients[1] = needle_read_chan.dmaClient;
   readClients[2] = mp_next_read_chan.dmaClient;

   Vector#(0, DMAWriteClient#(64)) writeClients = newVector();
`ifdef BSIM
   BsimDMAServer#(64) dma <- mkBsimDMAServer(dmaIndicationProxy.ifc, readClients, writeClients);
`else
   Integer numRequests = 8;
   AxiDMAServer#(64,8) dma <- mkAxiDMAServer(dmaIndicationProxy.ifc, numRequests, readClients, writeClients);
`endif
   DMARequestWrapper dmaRequestWrapper <- mkDMARequestWrapper(DMARequest,dma.request);

   StrstrIndicationProxy strstrIndicationProxy <- mkStrstrIndicationProxy(StrstrIndication);
   StrstrRequest strstrRequest <- mkStrstrRequest(strstrIndicationProxy.ifc, haystack_read_chan.dmaServer, 
						  needle_read_chan.dmaServer, mp_next_read_chan.dmaServer);
   StrstrRequestWrapper strstrRequestWrapper <- mkStrstrRequestWrapper(StrstrRequest,strstrRequest);

   Vector#(4,StdPortal) portals;
   portals[0] = strstrRequestWrapper.portalIfc;
   portals[1] = strstrIndicationProxy.portalIfc; 
   portals[2] = dmaRequestWrapper.portalIfc;
   portals[3] = dmaIndicationProxy.portalIfc; 
   
   Directory dir <- mkDirectory(portals);
   Vector#(1,StdPortal) directories;
   directories[0] = dir.portalIfc;
   
   // when constructing ctrl and interrupt muxes, directories must be the first argument
   let ctrl_mux <- mkAxiSlaveMux(directories,portals);
   let interrupt_mux <- mkInterruptMux(portals);
`ifndef BSIM
   let axi_master <- mkAxi3Master(dma.m_axi);
`endif
   
   interface ReadOnly interrupt = interrupt_mux;
   interface StdAxi3Slave ctrl = ctrl_mux;
`ifndef BSIM
   interface Vector m_axi = replicate(dma.m_axi);
`else
   interface Vector m_axi = ?;
`endif
   interface LEDS leds = ?;
endmodule
