// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;
import BRAM::*;
import DefaultValue::*;

// portz libraries
import Leds::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import PortalMemory::*;
import MemTypes::*;
import MemServer::*;

// generated by tool
import NandSimRequestWrapper::*;
import DmaConfigWrapper::*;
import StrstrRequestWrapper::*;

import NandSimIndicationProxy::*;
import DmaIndicationProxy::*;
import StrstrIndicationProxy::*;

// defined by user
import NandSim::*;
import Strstr::*;

typedef enum {DmaIndication, DmaConfig, NandSimIndication, NandSimRequest, StrstrIndication, StrstrRequest, StrstrDmaIndication, StrstrDmaConfig} IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalDmaTop#(PhysAddrWidth));
   
   NandSimIndicationProxy nandSimIndicationProxy <- mkNandSimIndicationProxy(NandSimIndication);
   NandSim#(1) nandSim <- mkNandSim(cons(nandSimIndicationProxy.ifc,nil));
   NandSimRequestWrapper nandSimRequestWrapper <- mkNandSimRequestWrapper(NandSimRequest,nandSim.requests[0]);
   
   StrstrIndicationProxy strstrIndicationProxy <- mkStrstrIndicationProxy(StrstrIndication);
   Strstr#(1,64) strstr <- mkStrstrRequest(strstrIndicationProxy.ifc);
   StrstrRequestWrapper strstrRequestWrapper <- mkStrstrRequestWrapper(StrstrRequest,strstr.request);

   DmaIndicationProxy dmaIndicationProxy <- mkDmaIndicationProxy(DmaIndication);
   MemServer#(PhysAddrWidth,64,1) dma <- mkMemServer(dmaIndicationProxy.ifc, cons(nandSim.readClient, nil), cons(nandSim.writeClient, nil));
   DmaConfigWrapper dmaRequestWrapper <- mkDmaConfigWrapper(DmaConfig,dma.request);
   
   DmaIndicationProxy strstrDmaIndicationProxy <- mkDmaIndicationProxy(StrstrDmaIndication);   
   MemServer#(PhysAddrWidth,64,1) strstrDma <- mkMemServerR(False, strstrDmaIndicationProxy.ifc, strstr.read_clients);
   DmaConfigWrapper strstrDmaRequestWrapper <- mkDmaConfigWrapper(StrstrDmaConfig, strstrDma.request);
   
   Vector#(8,StdPortal) portals;
   portals[0] = nandSimRequestWrapper.portalIfc;
   portals[1] = nandSimIndicationProxy.portalIfc; 
   portals[2] = dmaRequestWrapper.portalIfc;
   portals[3] = dmaIndicationProxy.portalIfc; 
   portals[4] = strstrRequestWrapper.portalIfc;
   portals[5] = strstrIndicationProxy.portalIfc; 
   portals[6] = strstrDmaRequestWrapper.portalIfc;
   portals[7] = strstrDmaIndicationProxy.portalIfc; 
   
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;
      
endmodule : mkPortalTop
