// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import AxiMasterSlave::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import BlueScope::*;
import PortalMemory::*;
import Dma::*;
import DmaUtils::*;
import PhysicalDma::*;

// generated by tool
import MaxcommonsubseqRequestWrapper::*;
import DmaConfigWrapper::*;
import MaxcommonsubseqIndicationProxy::*;
import DmaIndicationProxy::*;

// defined by user
import Maxcommonsubseq::*;

typedef enum {MaxcommonsubseqIndication, MaxcommonsubseqRequest, DmaIndication, DmaConfig} IfcNames deriving (Eq,Bits);
typedef 1 DegPar;


module mkPortalTop(StdPortalTop#(addrWidth)) 

   provisos(Add#(addrWidth, a__, 52),
	    Add#(b__, addrWidth, 64),
	    Add#(c__, 12, addrWidth),
	    Add#(addrWidth, d__, 44),
	    Add#(e__, c__, 40),
	    Add#(f__, addrWidth, 40));

   DmaIndicationProxy dmaIndicationProxy <- mkDmaIndicationProxy(DmaIndication);
   DmaReadBuffer#(64,1) setupA_read_chan <- mkDmaReadBuffer();
   DmaReadBuffer#(64,1) setupB_read_chan <- mkDmaReadBuffer();
   DmaWriteBuffer#(64,1) fetch_write_chan <- mkDmaWriteBuffer();
   
   DmaReadClient#(64) setupA_read_client = setupA_read_chan.dmaClient;
   DmaReadClient#(64) setupB_read_client = setupB_read_chan.dmaClient;
   DmaWriteClient#(64) fetch_write_client = fetch_write_chan.dmaClient;
   
   Vector#(2,  DmaReadClient#(64)) readClients;
   readClients[0] = setupA_read_client;
   readClients[1] = setupB_read_client;

   Vector#(1, DmaWriteClient#(64)) writeClients;
   writeClients[0] = fetch_write_client;


   PhysicalDmaServer#(addrWidth,64) dma <- mkPhysicalDmaServer(dmaIndicationProxy.ifc, readClients, writeClients);
   
   DmaConfigWrapper dmaConfigWrapper <- mkDmaConfigWrapper(DmaConfig, dma.request);
   
   MaxcommonsubseqIndicationProxy maxcommonsubseqIndicationProxy <- mkMaxcommonsubseqIndicationProxy(MaxcommonsubseqIndication);
   MaxcommonsubseqRequest maxcommonsubseqRequest <- mkMaxcommonsubseqRequest(maxcommonsubseqIndicationProxy.ifc, setupA_read_chan.dmaServer, setupB_read_chan.dmaServer, fetch_write_chan.dmaServer);
   MaxcommonsubseqRequestWrapper maxcommonsubseqRequestWrapper <- mkMaxcommonsubseqRequestWrapper(MaxcommonsubseqRequest,maxcommonsubseqRequest);

   Vector#(4,StdPortal) portals;
   portals[0] = maxcommonsubseqRequestWrapper.portalIfc;
   portals[1] = maxcommonsubseqIndicationProxy.portalIfc; 
   portals[2] = dmaConfigWrapper.portalIfc;
   portals[3] = dmaIndicationProxy.portalIfc; 
   
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkAxiSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface ctrl = ctrl_mux;
   interface read_client = dma.read_client;
   interface write_client = dma.write_client;
   interface leds = default_leds;
endmodule
