// bsv libraries
import Vector::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import MemTypes::*;
import MemPortal::*;

// generated by tool
import Tiny3IndicationProxy::*;
import Tiny3RequestWrapper::*;

// defined by user
import Tiny3::*;

typedef enum {Tiny3Indication, Tiny3Request} IfcNames deriving (Eq,Bits);

module mkConnectalTop(StdConnectalTop#(PhysAddrWidth));

   // instantiate user portals
   Tiny3IndicationProxy tiny3IndicationProxy <- mkTiny3IndicationProxy(Tiny3Indication);
   Tiny3Request tiny3Request <- mkTiny3Request(tiny3IndicationProxy.ifc);
   Tiny3RequestWrapper tiny3RequestWrapper <- mkTiny3RequestWrapper(Tiny3Request,tiny3Request);
   
   Vector#(2,StdPortal) portals;
   portals[0] = tiny3RequestWrapper.portalIfc;
   portals[1] = tiny3IndicationProxy.portalIfc;
   
   // instantiate system directory
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = nil;
   interface leds = default_leds;

endmodule : mkConnectalTop


