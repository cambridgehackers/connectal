// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import CtrlMux::*;
import Portal::*;
import Leds::*;
import ConnectalMemory::*;
import MemServer::*;
import MMU::*;
import ConnectalMemory::*;
import MemTypes::*;
import MemUtils::*;
import RbmTypes::*;
import HostInterface::*;

// generated by tool
import DmaDebugRequest::*;
import MMUConfigRequest::*;
import DmaDebugIndication::*;
import MMUConfigIndication::*;

module  mkConnectalTop#(HostType host)(ConnectalTop#(PhysAddrWidth,TMul#(32,N),Empty,NumberOfMasters));

   // all this stuff is here so we can call portalAlloc in user space
   let reader <- mkMemReader();
   let writer <- mkMemWriter();

   Vector#(1,MemReadClient#(TMul#(32,N)))  readClients  = cons(reader.readClient, nil);
   Vector#(1,MemWriteClient#(TMul#(32,N))) writeClients = cons(writer.writeClient, nil);

   MMUConfigIndicationProxy hostMMUConfigIndicationProxy <- mkMMUConfigIndicationProxy(HostMMUConfigIndication);
   MMU#(PhysAddrWidth) hostMMU <- mkMMU(0, True, hostMMUConfigIndicationProxy.ifc);
   MMUConfigRequestWrapper hostMMUConfigRequestWrapper <- mkMMUConfigRequestWrapper(HostMMUConfigRequest, hostMMU.request);

   DmaDebugIndicationProxy hostDmaDebugIndicationProxy <- mkDmaDebugIndicationProxy(HostDmaDebugIndication);
   MemServer#(PhysAddrWidth,TMul#(32,N), NumberOfMasters) dma <- mkMemServerRW(hostMMUConfigIndicationProxy.ifc,
									       hostDmaDebugIndicationProxy.ifc, readClients, writeClients, cons(hostMMU,nil));
   DmaDebugRequestWrapper hostDmaDebugRequestWrapper <- mkDmaDebugRequestWrapper(HostDmaDebugRequest, dma.request);

   Vector#(4,StdPortal) portals;
   portals[0] = hostDmaDebugIndicationProxy.portalIfc; 
   portals[1] = hostDmaDebugRequestWrapper.portalIfc;
   portals[2] = hostMMUConfigRequestWrapper.portalIfc;
   portals[3] = hostMMUConfigIndicationProxy.portalIfc;
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;

endmodule : mkConnectalTop
