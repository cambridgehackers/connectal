// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import PortalMemory::*;
import MemTypes::*;
import MemServer::*;

// generated by tool
import GrepRequestWrapper::*;
import DmaConfigWrapper::*;
import GrepIndicationProxy::*;
import DmaIndicationProxy::*;

// defined by user
import Grep::*;

typedef enum {GrepIndication, GrepRequest, DmaIndication, DmaConfig} IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalDmaTop#(PhysAddrWidth));

   GrepIndicationProxy grepIndicationProxy <- mkGrepIndicationProxy(GrepIndication);
   Grep#(64) grep <- mkGrep(grepIndicationProxy.ifc);
   GrepRequestWrapper grepRequestWrapper <- mkGrepRequestWrapper(GrepRequest,grep.request);
   
   let read_clients = cons(grep.config_read_client, cons(grep.haystack_read_client,nil));
   DmaIndicationProxy dmaIndicationProxy <- mkDmaIndicationProxy(DmaIndication);
   MemServer#(PhysAddrWidth,64,1) dma <- mkMemServerR(True, dmaIndicationProxy.ifc, read_clients);
   DmaConfigWrapper dmaConfigWrapper <- mkDmaConfigWrapper(DmaConfig, dma.request);

   Vector#(4,StdPortal) portals;
   portals[0] = grepRequestWrapper.portalIfc;
   portals[1] = grepIndicationProxy.portalIfc; 
   portals[2] = dmaConfigWrapper.portalIfc;
   portals[3] = dmaIndicationProxy.portalIfc; 
   
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;
endmodule
