// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;

// portz libraries
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import BlueScope::*;
import PortalMemory::*;
import MemTypes::*;
import DmaUtils::*;
import MemServer::*;

// generated by tool
import SpliceRequestWrapper::*;
import DmaConfigWrapper::*;
import SpliceIndicationProxy::*;
import DmaIndicationProxy::*;

// defined by user
import Splice::*;

typedef enum {SpliceIndication, SpliceRequest, DmaIndication, DmaConfig} IfcNames deriving (Eq,Bits);
typedef 1 DegPar;


module mkPortalTop(StdPortalDmaTop#(addrWidth)) 

   provisos(Add#(addrWidth, a__, 52),
	    Add#(b__, addrWidth, 64),
	    Add#(c__, 12, addrWidth),
	    Add#(addrWidth, d__, 44),
	    Add#(e__, c__, 40),
	    Add#(f__, addrWidth, 40));

   DmaIndicationProxy dmaIndicationProxy <- mkDmaIndicationProxy(DmaIndication);
   DmaReadBuffer#(64,1) setupA_read_chan <- mkDmaReadBuffer();
   DmaReadBuffer#(64,1) setupB_read_chan <- mkDmaReadBuffer();
   DmaWriteBuffer#(64,1) fetch_write_chan <- mkDmaWriteBuffer();
   
   ObjectReadClient#(64) setupA_read_client = setupA_read_chan.dmaClient;
   ObjectReadClient#(64) setupB_read_client = setupB_read_chan.dmaClient;
   ObjectWriteClient#(64) fetch_write_client = fetch_write_chan.dmaClient;
   
   Vector#(2,  ObjectReadClient#(64)) readClients;
   readClients[0] = setupA_read_client;
   readClients[1] = setupB_read_client;

   Vector#(1, ObjectWriteClient#(64)) writeClients;
   writeClients[0] = fetch_write_client;


   MemServer#(addrWidth,64,1) dma <- mkMemServer(dmaIndicationProxy.ifc, readClients, writeClients);
   
   DmaConfigWrapper dmaConfigWrapper <- mkDmaConfigWrapper(DmaConfig, dma.request);
   
   SpliceIndicationProxy spliceIndicationProxy <- mkSpliceIndicationProxy(SpliceIndication);
   SpliceRequest spliceRequest <- mkSpliceRequest(spliceIndicationProxy.ifc, setupA_read_chan.dmaServer, setupB_read_chan.dmaServer, fetch_write_chan.dmaServer);
   SpliceRequestWrapper spliceRequestWrapper <- mkSpliceRequestWrapper(SpliceRequest,spliceRequest);

   Vector#(4,StdPortal) portals;
   portals[0] = spliceRequestWrapper.portalIfc;
   portals[1] = spliceIndicationProxy.portalIfc; 
   portals[2] = dmaConfigWrapper.portalIfc;
   portals[3] = dmaIndicationProxy.portalIfc; 
   
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;
endmodule
