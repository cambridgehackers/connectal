
module axi_passthrough ();
endmodule
