// Copyright (c) 2013 Nokia, Inc.
// Copyright (c) 2013 Quanta Research Cambridge, Inc.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.
import Clocks::*;
import FIFO::*;
import GetPut::*;
import Vector::*;

interface EchoIndication;
    method Action heard(Bit#(32) v);
    method Action heard2(Bit#(16) a, Bit#(16) b);
endinterface

interface EchoRequest;
   method Action say(Bit#(32) v);
   method Action say2(Bit#(16) a, Bit#(16) b);
   method Action setLeds(Bit#(8) v);
endinterface

interface Echo;
   interface EchoRequest request;
endinterface

typedef struct {
	Bit#(16) a;
	Bit#(16) b;
} EchoPair deriving (Bits);

module mkEcho#(Clock derivedClock, Reset derivedReset, EchoIndication indication)(Echo);
   let clock <- exposeCurrentClock;
   let reset <- exposeCurrentReset;

    let delay_toslow <- mkSyncFIFO(16, clock, reset, derivedClock);
    let delay_fromslow <- mkSyncFIFO(16, derivedClock, derivedReset, clock);
    let delay2_toslow <- mkSyncFIFO(16, clock, reset, derivedClock);
    let delay2_fromslow <- mkSyncFIFO(16, derivedClock, derivedReset, clock);

   rule heard_slow; // derivedClock domain
      let v <- toGet(delay_toslow).get();
      delay_fromslow.enq(v);
   endrule
   rule hear_fast;
      let v <- toGet(delay_fromslow).get();
      indication.heard(v);
   endrule

   rule heard2_slow; // derivedClock domain
      let v <- toGet(delay2_toslow).get();
      delay2_fromslow.enq(v);
   endrule
   rule heard2_fast;
      let v <- toGet(delay2_fromslow).get();
      indication.heard2(v.b, v.a);
   endrule
   
   interface EchoRequest request;
      method Action say(Bit#(32) v);
	 delay_toslow.enq(v);
      endmethod
      
      method Action say2(Bit#(16) a, Bit#(16) b);
	 delay2_toslow.enq(EchoPair { a: a, b: b});
      endmethod
      
      method Action setLeds(Bit#(8) v);
      endmethod
   endinterface
endmodule
