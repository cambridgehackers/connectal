// bsv libraries
import Vector::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import Portal::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import AxiMasterSlave::*;

// generated by tool
import SinkIndicationProxy::*;
import SinkRequestWrapper::*;

// defined by user
import Sink::*;

typedef enum {SinkIndication, SinkRequest} IfcNames deriving (Eq,Bits);

module mkPortalTop(StdPortalTop#(addrWidth));

   // instantiate user portals
   SinkIndicationProxy sinkIndicationProxy <- mkSinkIndicationProxy(SinkIndication);
   SinkRequest sinkRequest <- mkSinkRequest(sinkIndicationProxy.ifc);
   SinkRequestWrapper sinkRequestWrapper <- mkSinkRequestWrapper(SinkRequest,sinkRequest);
   
   Vector#(2,StdPortal) portals;
   portals[0] = sinkIndicationProxy.portalIfc;
   portals[1] = sinkRequestWrapper.portalIfc; 
   
   // instantiate system directory
   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkAxiSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface ctrl = ctrl_mux;
   interface m_axi = null_axi_master;
   interface leds = default_leds;

endmodule : mkPortalTop
