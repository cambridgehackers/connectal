
import Clocks::*;
import DefaultValue::*;
import XilinxCells::*;
import GetPut::*;

interface Pps7Can#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      phy_rx(Bit#(1) v);
    method Bit#(1)     phy_tx();
endinterface
interface Pps7Core#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      nfiq(Bit#(1) v);
    method Action      nirq(Bit#(1) v);
endinterface
interface Pps7Ddr#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      arb(Bit#(4) v);
    interface Inout#(Bit#(15))     addr;
    interface Inout#(Bit#(3))     bankaddr;
    interface Inout#(Bit#(1))     cas_n;
    interface Inout#(Bit#(1))     cke;
    interface Inout#(Bit#(1))     cs_n;
    interface Inout#(Bit#(1))     clk;
    interface Inout#(Bit#(1))     clk_n;
    interface Inout#(Bit#(c_dm_width))     dm;
    interface Inout#(Bit#(c_dq_width))     dq;
    interface Inout#(Bit#(c_dqs_width))     dqs;
    interface Inout#(Bit#(c_dqs_width))     dqs_n;
    interface Inout#(Bit#(1))     drstb;
    interface Inout#(Bit#(1))     odt;
    interface Inout#(Bit#(1))     ras_n;
    interface Inout#(Bit#(1))     vrn;
    interface Inout#(Bit#(1))     vrp;
    interface Inout#(Bit#(1))     web;
endinterface
interface Pps7Dma#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      aclk(Bit#(1) v);
    method Action      daready(Bit#(1) v);
    method Bit#(2)     datype();
    method Bit#(1)     davalid();
    method Action      drlast(Bit#(1) v);
    method Bit#(1)     drready();
    method Action      drtype(Bit#(2) v);
    method Action      drvalid(Bit#(1) v);
    method Bit#(1)     rstn();
endinterface
interface Pps7Enet#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      ext_intin(Bit#(1) v);
    method Action      gmii_col(Bit#(1) v);
    method Action      gmii_crs(Bit#(1) v);
    method Action      gmii_rxd(Bit#(8) v);
    method Action      gmii_rx_clk(Bit#(1) v);
    method Action      gmii_rx_dv(Bit#(1) v);
    method Action      gmii_rx_er(Bit#(1) v);
    method Bit#(8)     gmii_txd();
    method Action      gmii_tx_clk(Bit#(1) v);
    method Bit#(1)     gmii_tx_en();
    method Bit#(1)     gmii_tx_er();
    method Action      mdio_i(Bit#(1) v);
    method Bit#(1)     mdio_mdc();
    method Bit#(1)     mdio_o();
    method Bit#(1)     mdio_t();
    method Bit#(1)     ptp_delay_req_rx();
    method Bit#(1)     ptp_delay_req_tx();
    method Bit#(1)     ptp_pdelay_req_rx();
    method Bit#(1)     ptp_pdelay_req_tx();
    method Bit#(1)     ptp_pdelay_resp_rx();
    method Bit#(1)     ptp_pdelay_resp_tx();
    method Bit#(1)     ptp_sync_frame_rx();
    method Bit#(1)     ptp_sync_frame_tx();
    method Bit#(1)     sof_rx();
    method Bit#(1)     sof_tx();
endinterface
interface Pps7Event#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      eventi(Bit#(1) v);
    method Bit#(1)     evento();
    method Bit#(2)     standbywfe();
    method Bit#(2)     standbywfi();
endinterface
interface Pps7Fclk#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Bit#(1)     clk0();
    method Bit#(1)     clk1();
    method Bit#(1)     clk2();
    method Bit#(1)     clk3();
endinterface
interface Pps7Fclk_clktrig#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      n(Bit#(1) v);
endinterface
interface Pps7Fclk_reset#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Bit#(1)     n();
endinterface
interface Pps7Fpga#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      idle_n(Bit#(1) v);
endinterface
interface Pps7Ftmd#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      tracein_atid(Bit#(4) v);
    method Action      tracein_clk(Bit#(1) v);
    method Action      tracein_data(Bit#(32) v);
    method Action      tracein_valid(Bit#(1) v);
endinterface
interface Pps7Ftmt#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      f2p_debug(Bit#(32) v);
    method Action      f2p_trig(Bit#(4) v);
    method Bit#(4)     f2p_trigack();
    method Bit#(32)     p2f_debug();
    method Bit#(4)     p2f_trig();
    method Action      p2f_trigack(Bit#(4) v);
endinterface
interface Pps7Gpio#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      i(Bit#(gpio_width) v);
    method Bit#(gpio_width)     o();
    method Bit#(gpio_width)     t();
endinterface
interface Pps7I2c#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      scl_i(Bit#(1) v);
    method Bit#(1)     scl_o();
    method Bit#(1)     scl_t();
    method Action      sda_i(Bit#(1) v);
    method Bit#(1)     sda_o();
    method Bit#(1)     sda_t();
endinterface
interface Pps7Irq#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      f2p(Bit#(16) v);
    method Bit#(1)     p2f_can0();
    method Bit#(1)     p2f_can1();
    method Bit#(1)     p2f_cti();
    method Bit#(1)     p2f_dmac0();
    method Bit#(1)     p2f_dmac1();
    method Bit#(1)     p2f_dmac2();
    method Bit#(1)     p2f_dmac3();
    method Bit#(1)     p2f_dmac4();
    method Bit#(1)     p2f_dmac5();
    method Bit#(1)     p2f_dmac6();
    method Bit#(1)     p2f_dmac7();
    method Bit#(1)     p2f_dmac_abort();
    method Bit#(1)     p2f_enet0();
    method Bit#(1)     p2f_enet1();
    method Bit#(1)     p2f_enet_wake0();
    method Bit#(1)     p2f_enet_wake1();
    method Bit#(1)     p2f_gpio();
    method Bit#(1)     p2f_i2c0();
    method Bit#(1)     p2f_i2c1();
    method Bit#(1)     p2f_qspi();
    method Bit#(1)     p2f_sdio0();
    method Bit#(1)     p2f_sdio1();
    method Bit#(1)     p2f_smc();
    method Bit#(1)     p2f_spi0();
    method Bit#(1)     p2f_spi1();
    method Bit#(1)     p2f_uart0();
    method Bit#(1)     p2f_uart1();
    method Bit#(1)     p2f_usb0();
    method Bit#(1)     p2f_usb1();
endinterface
interface Pps7M_axi_gp#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      aclk(Bit#(1) v);
    method Bit#(32)     araddr();
    method Bit#(2)     arburst();
    method Bit#(4)     arcache();
    method Bit#(1)     aresetn();
    method Bit#(id_width)     arid();
    method Bit#(4)     arlen();
    method Bit#(2)     arlock();
    method Bit#(3)     arprot();
    method Bit#(4)     arqos();
    method Action      arready(Bit#(1) v);
    method Bit#(3)     arsize();
    method Bit#(1)     arvalid();
    method Bit#(32)     awaddr();
    method Bit#(2)     awburst();
    method Bit#(4)     awcache();
    method Bit#(id_width)     awid();
    method Bit#(4)     awlen();
    method Bit#(2)     awlock();
    method Bit#(3)     awprot();
    method Bit#(4)     awqos();
    method Action      awready(Bit#(1) v);
    method Bit#(3)     awsize();
    method Bit#(1)     awvalid();
    method Action      bid(Bit#(id_width) v);
    method Bit#(1)     bready();
    method Action      bresp(Bit#(2) v);
    method Action      bvalid(Bit#(1) v);
    method Action      rdata(Bit#(32) v);
    method Action      rid(Bit#(id_width) v);
    method Action      rlast(Bit#(1) v);
    method Bit#(1)     rready();
    method Action      rresp(Bit#(2) v);
    method Action      rvalid(Bit#(1) v);
    method Bit#(32)     wdata();
    method Bit#(id_width)     wid();
    method Bit#(1)     wlast();
    method Action      wready(Bit#(1) v);
    method Bit#(4)     wstrb();
    method Bit#(1)     wvalid();
endinterface
interface Pps7Pjtag#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      tck(Bit#(1) v);
    method Action      td_i(Bit#(1) v);
    method Bit#(1)     td_o();
    method Bit#(1)     td_t();
    method Action      tms(Bit#(1) v);
endinterface
interface Pps7Ps#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      clk(Bit#(1) v);
    method Action      porb(Bit#(1) v);
    method Action      srstb(Bit#(1) v);
endinterface
interface Pps7S_axi_acp#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      aclk(Bit#(1) v);
    method Action      araddr(Bit#(32) v);
    method Action      arburst(Bit#(2) v);
    method Action      arcache(Bit#(4) v);
    method Bit#(1)     aresetn();
    method Action      arid(Bit#(id_width) v);
    method Action      arlen(Bit#(4) v);
    method Action      arlock(Bit#(2) v);
    method Action      arprot(Bit#(3) v);
    method Action      arqos(Bit#(4) v);
    method Bit#(1)     arready();
    method Action      arsize(Bit#(3) v);
    method Action      aruser(Bit#(5) v);
    method Action      arvalid(Bit#(1) v);
    method Action      awaddr(Bit#(32) v);
    method Action      awburst(Bit#(2) v);
    method Action      awcache(Bit#(4) v);
    method Action      awid(Bit#(id_width) v);
    method Action      awlen(Bit#(4) v);
    method Action      awlock(Bit#(2) v);
    method Action      awprot(Bit#(3) v);
    method Action      awqos(Bit#(4) v);
    method Bit#(1)     awready();
    method Action      awsize(Bit#(3) v);
    method Action      awuser(Bit#(5) v);
    method Action      awvalid(Bit#(1) v);
    method Bit#(id_width)     bid();
    method Action      bready(Bit#(1) v);
    method Bit#(2)     bresp();
    method Bit#(1)     bvalid();
    method Bit#(64)     rdata();
    method Bit#(id_width)     rid();
    method Bit#(1)     rlast();
    method Action      rready(Bit#(1) v);
    method Bit#(2)     rresp();
    method Bit#(1)     rvalid();
    method Action      wdata(Bit#(64) v);
    method Action      wid(Bit#(id_width) v);
    method Action      wlast(Bit#(1) v);
    method Bit#(1)     wready();
    method Action      wstrb(Bit#(8) v);
    method Action      wvalid(Bit#(1) v);
endinterface
interface Pps7S_axi_gp#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      aclk(Bit#(1) v);
    method Action      araddr(Bit#(32) v);
    method Action      arburst(Bit#(2) v);
    method Action      arcache(Bit#(4) v);
    method Bit#(1)     aresetn();
    method Action      arid(Bit#(id_width) v);
    method Action      arlen(Bit#(4) v);
    method Action      arlock(Bit#(2) v);
    method Action      arprot(Bit#(3) v);
    method Action      arqos(Bit#(4) v);
    method Bit#(1)     arready();
    method Action      arsize(Bit#(3) v);
    method Action      arvalid(Bit#(1) v);
    method Action      awaddr(Bit#(32) v);
    method Action      awburst(Bit#(2) v);
    method Action      awcache(Bit#(4) v);
    method Action      awid(Bit#(id_width) v);
    method Action      awlen(Bit#(4) v);
    method Action      awlock(Bit#(2) v);
    method Action      awprot(Bit#(3) v);
    method Action      awqos(Bit#(4) v);
    method Bit#(1)     awready();
    method Action      awsize(Bit#(3) v);
    method Action      awvalid(Bit#(1) v);
    method Bit#(id_width)     bid();
    method Action      bready(Bit#(1) v);
    method Bit#(2)     bresp();
    method Bit#(1)     bvalid();
    method Bit#(32)     rdata();
    method Bit#(id_width)     rid();
    method Bit#(1)     rlast();
    method Action      rready(Bit#(1) v);
    method Bit#(2)     rresp();
    method Bit#(1)     rvalid();
    method Action      wdata(Bit#(32) v);
    method Action      wid(Bit#(id_width) v);
    method Action      wlast(Bit#(1) v);
    method Bit#(1)     wready();
    method Action      wstrb(Bit#(4) v);
    method Action      wvalid(Bit#(1) v);
endinterface
interface Pps7S_axi_hp#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      aclk(Bit#(1) v);
    method Action      araddr(Bit#(32) v);
    method Action      arburst(Bit#(2) v);
    method Action      arcache(Bit#(4) v);
    method Bit#(1)     aresetn();
    method Action      arid(Bit#(id_width) v);
    method Action      arlen(Bit#(4) v);
    method Action      arlock(Bit#(2) v);
    method Action      arprot(Bit#(3) v);
    method Action      arqos(Bit#(4) v);
    method Bit#(1)     arready();
    method Action      arsize(Bit#(3) v);
    method Action      arvalid(Bit#(1) v);
    method Action      awaddr(Bit#(32) v);
    method Action      awburst(Bit#(2) v);
    method Action      awcache(Bit#(4) v);
    method Action      awid(Bit#(id_width) v);
    method Action      awlen(Bit#(4) v);
    method Action      awlock(Bit#(2) v);
    method Action      awprot(Bit#(3) v);
    method Action      awqos(Bit#(4) v);
    method Bit#(1)     awready();
    method Action      awsize(Bit#(3) v);
    method Action      awvalid(Bit#(1) v);
    method Bit#(id_width)     bid();
    method Action      bready(Bit#(1) v);
    method Bit#(2)     bresp();
    method Bit#(1)     bvalid();
    method Bit#(3)     racount();
    method Bit#(8)     rcount();
    method Bit#(data_width)     rdata();
    method Action      rdissuecap1_en(Bit#(1) v);
    method Bit#(id_width)     rid();
    method Bit#(1)     rlast();
    method Action      rready(Bit#(1) v);
    method Bit#(2)     rresp();
    method Bit#(1)     rvalid();
    method Bit#(6)     wacount();
    method Bit#(8)     wcount();
    method Action      wdata(Bit#(data_width) v);
    method Action      wid(Bit#(id_width) v);
    method Action      wlast(Bit#(1) v);
    method Bit#(1)     wready();
    method Action      wrissuecap1_en(Bit#(1) v);
    method Action      wstrb(Bit#(TDiv#(data_width,8)) v);
    method Action      wvalid(Bit#(1) v);
endinterface
interface Pps7Sdio#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Bit#(1)     buspow();
    method Bit#(3)     busvolt();
    method Action      cdn(Bit#(1) v);
    method Bit#(1)     clk();
    method Action      clk_fb(Bit#(1) v);
    method Action      cmd_i(Bit#(1) v);
    method Bit#(1)     cmd_o();
    method Bit#(1)     cmd_t();
    method Action      data_i(Bit#(4) v);
    method Bit#(4)     data_o();
    method Bit#(4)     data_t();
    method Bit#(1)     led();
    method Action      wp(Bit#(1) v);
endinterface
interface Pps7Spi#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      miso_i(Bit#(1) v);
    method Bit#(1)     miso_o();
    method Bit#(1)     miso_t();
    method Action      mosi_i(Bit#(1) v);
    method Bit#(1)     mosi_o();
    method Bit#(1)     mosi_t();
    method Action      sclk_i(Bit#(1) v);
    method Bit#(1)     sclk_o();
    method Bit#(1)     sclk_t();
    method Bit#(1)     ss1_o();
    method Bit#(1)     ss2_o();
    method Action      ss_i(Bit#(1) v);
    method Bit#(1)     ss_o();
    method Bit#(1)     ss_t();
endinterface
interface Pps7Sram#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      intin(Bit#(1) v);
endinterface
interface Pps7Trace#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      clk(Bit#(1) v);
    method Bit#(1)     ctl();
    method Bit#(32)     data();
endinterface
interface Pps7Ttc#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      clk0_in(Bit#(1) v);
    method Action      clk1_in(Bit#(1) v);
    method Action      clk2_in(Bit#(1) v);
    method Bit#(1)     wave0_out();
    method Bit#(1)     wave1_out();
    method Bit#(1)     wave2_out();
endinterface
interface Pps7Uart#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      ctsn(Bit#(1) v);
    method Action      dcdn(Bit#(1) v);
    method Action      dsrn(Bit#(1) v);
    method Bit#(1)     dtrn();
    method Action      rin(Bit#(1) v);
    method Bit#(1)     rtsn();
    method Action      rx(Bit#(1) v);
    method Bit#(1)     tx();
endinterface
interface Pps7Usb#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Bit#(2)     port_indctl();
    method Action      vbus_pwrfault(Bit#(1) v);
    method Bit#(1)     vbus_pwrselect();
endinterface
interface Pps7Wdt#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    method Action      clk_in(Bit#(1) v);
    method Bit#(1)     rst_out();
endinterface
interface PPS7#(numeric type c_dm_width, numeric type c_dq_width, numeric type c_dqs_width, numeric type data_width, numeric type gpio_width, numeric type id_width, numeric type mio_width);
    interface Pps7Can#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     can0;
    interface Pps7Can#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     can1;
    interface Pps7Core#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     core0;
    interface Pps7Core#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     core1;
    interface Pps7Ddr#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     ddr;
    interface Pps7Dma#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     dma0;
    interface Pps7Dma#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     dma1;
    interface Pps7Dma#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     dma2;
    interface Pps7Dma#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     dma3;
    interface Pps7Enet#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     enet0;
    interface Pps7Enet#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     enet1;
    interface Pps7Event#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     event_;
    interface Pps7Fclk#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     fclk;
    interface Pps7Fclk_clktrig#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     fclk_clktrig0;
    interface Pps7Fclk_clktrig#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     fclk_clktrig1;
    interface Pps7Fclk_clktrig#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     fclk_clktrig2;
    interface Pps7Fclk_clktrig#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     fclk_clktrig3;
    interface Pps7Fclk_reset#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     fclk_reset0;
    interface Pps7Fclk_reset#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     fclk_reset1;
    interface Pps7Fclk_reset#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     fclk_reset2;
    interface Pps7Fclk_reset#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     fclk_reset3;
    interface Pps7Fpga#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     fpga;
    interface Pps7Ftmd#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     ftmd;
    interface Pps7Ftmt#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     ftmt;
    interface Pps7Gpio#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     gpio;
    interface Pps7I2c#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     i2c0;
    interface Pps7I2c#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     i2c1;
    interface Pps7Irq#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     irq;
    interface Inout#(Bit#(mio_width))     mio;
    interface Pps7M_axi_gp#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     m_axi_gp0;
    interface Pps7M_axi_gp#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     m_axi_gp1;
    interface Pps7Pjtag#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     pjtag;
    interface Pps7Ps#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     ps;
    interface Pps7Sdio#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     sdio0;
    interface Pps7Sdio#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     sdio1;
    interface Pps7Spi#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     spi0;
    interface Pps7Spi#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     spi1;
    interface Pps7Sram#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     sram;
    interface Pps7S_axi_acp#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     s_axi_acp;
    interface Pps7S_axi_gp#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     s_axi_gp0;
    interface Pps7S_axi_gp#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     s_axi_gp1;
    interface Pps7S_axi_hp#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     s_axi_hp0;
    interface Pps7S_axi_hp#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     s_axi_hp1;
    interface Pps7S_axi_hp#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     s_axi_hp2;
    interface Pps7S_axi_hp#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     s_axi_hp3;
    interface Pps7Trace#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     trace;
    interface Pps7Ttc#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     ttc0;
    interface Pps7Ttc#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     ttc1;
    interface Pps7Uart#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     uart0;
    interface Pps7Uart#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     uart1;
    interface Pps7Usb#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     usb0;
    interface Pps7Usb#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     usb1;
    interface Pps7Wdt#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width)     wdt;
endinterface
import "BVI" processing_system7 =
module mkPPS7(PPS7#(c_dm_width, c_dq_width, c_dqs_width, data_width, gpio_width, id_width, mio_width));
    let c_dm_width = valueOf(c_dm_width);
    let c_dq_width = valueOf(c_dq_width);
    let c_dqs_width = valueOf(c_dqs_width);
    let data_width = valueOf(data_width);
    let gpio_width = valueOf(gpio_width);
    let id_width = valueOf(id_width);
    let mio_width = valueOf(mio_width);
    parameter C_DM_WIDTH = 4;
    parameter C_DQS_WIDTH = 4;
    parameter C_DQ_WIDTH = 32;
    parameter C_EMIO_GPIO_WIDTH = 64;
    parameter C_EN_EMIO_ENET0 = 0;
    parameter C_EN_EMIO_ENET1 = 0;
    parameter C_EN_EMIO_TRACE = 0;
    parameter C_FCLK_CLK0_BUF = "TRUE";
    parameter C_FCLK_CLK1_BUF = "TRUE";
    parameter C_FCLK_CLK2_BUF = "TRUE";
    parameter C_FCLK_CLK3_BUF = "TRUE";
    parameter C_INCLUDE_ACP_TRANS_CHECK = 0;
    parameter C_INCLUDE_TRACE_BUFFER = 0;
    parameter C_MIO_PRIMITIVE = 54;
    parameter C_M_AXI_GP0_ENABLE_STATIC_REMAP = 1;
    parameter C_M_AXI_GP0_ID_WIDTH = 12;
    parameter C_M_AXI_GP0_THREAD_ID_WIDTH = 12;
    parameter C_M_AXI_GP1_ENABLE_STATIC_REMAP = 1;
    parameter C_M_AXI_GP1_ID_WIDTH = 12;
    parameter C_M_AXI_GP1_THREAD_ID_WIDTH = 12;
    parameter C_NUM_F2P_INTR_INPUTS = 2;
    parameter C_PACKAGE_NAME = "clg484";
    parameter C_PS7_SI_REV = "PRODUCTION";
    parameter C_S_AXI_ACP_ARUSER_VAL = 31;
    parameter C_S_AXI_ACP_AWUSER_VAL = 31;
    parameter C_S_AXI_ACP_ID_WIDTH = 3;
    parameter C_S_AXI_GP0_ID_WIDTH = 6;
    parameter C_S_AXI_GP1_ID_WIDTH = 6;
    parameter C_S_AXI_HP0_DATA_WIDTH = 64;
    parameter C_S_AXI_HP0_ID_WIDTH = 6;
    parameter C_S_AXI_HP1_DATA_WIDTH = 64;
    parameter C_S_AXI_HP1_ID_WIDTH = 6;
    parameter C_S_AXI_HP2_DATA_WIDTH = 64;
    parameter C_S_AXI_HP2_ID_WIDTH = 6;
    parameter C_S_AXI_HP3_DATA_WIDTH = 64;
    parameter C_S_AXI_HP3_ID_WIDTH = 6;
    parameter C_TRACE_BUFFER_CLOCK_DELAY = 12;
    parameter C_TRACE_BUFFER_FIFO_SIZE = 128;
    parameter C_USE_DEFAULT_ACP_USER_VAL = 1;
    parameter USE_TRACE_DATA_EDGE_DETECTOR = 0;
    interface Pps7Can     can0;
        method phy_rx(CAN0_PHY_RX) enable((*inhigh*) en100);
        method CAN0_PHY_TX phy_tx();
    endinterface
    interface Pps7Can     can1;
        method phy_rx(CAN1_PHY_RX) enable((*inhigh*) en101);
        method CAN1_PHY_TX phy_tx();
    endinterface
    interface Pps7Core     core0;
        method nfiq(Core0_nFIQ) enable((*inhigh*) en102);
        method nirq(Core0_nIRQ) enable((*inhigh*) en103);
    endinterface
    interface Pps7Core     core1;
        method nfiq(Core1_nFIQ) enable((*inhigh*) en104);
        method nirq(Core1_nIRQ) enable((*inhigh*) en105);
    endinterface
    interface Pps7Ddr     ddr;
        method arb(DDR_ARB) enable((*inhigh*) en106);
        ifc_inout addr(DDR_Addr);
        ifc_inout bankaddr(DDR_BankAddr);
        ifc_inout cas_n(DDR_CAS_n);
        ifc_inout cke(DDR_CKE);
        ifc_inout cs_n(DDR_CS_n);
        ifc_inout clk(DDR_Clk);
        ifc_inout clk_n(DDR_Clk_n);
        ifc_inout dm(DDR_DM);
        ifc_inout dq(DDR_DQ);
        ifc_inout dqs(DDR_DQS);
        ifc_inout dqs_n(DDR_DQS_n);
        ifc_inout drstb(DDR_DRSTB);
        ifc_inout odt(DDR_ODT);
        ifc_inout ras_n(DDR_RAS_n);
        ifc_inout vrn(DDR_VRN);
        ifc_inout vrp(DDR_VRP);
        ifc_inout web(DDR_WEB);
    endinterface
    interface Pps7Dma     dma0;
        method aclk(DMA0_ACLK) enable((*inhigh*) en107);
        method daready(DMA0_DAREADY) enable((*inhigh*) en108);
        method DMA0_DATYPE datype();
        method DMA0_DAVALID davalid();
        method drlast(DMA0_DRLAST) enable((*inhigh*) en109);
        method DMA0_DRREADY drready();
        method drtype(DMA0_DRTYPE) enable((*inhigh*) en110);
        method drvalid(DMA0_DRVALID) enable((*inhigh*) en111);
        method DMA0_RSTN rstn();
    endinterface
    interface Pps7Dma     dma1;
        method aclk(DMA1_ACLK) enable((*inhigh*) en112);
        method daready(DMA1_DAREADY) enable((*inhigh*) en113);
        method DMA1_DATYPE datype();
        method DMA1_DAVALID davalid();
        method drlast(DMA1_DRLAST) enable((*inhigh*) en114);
        method DMA1_DRREADY drready();
        method drtype(DMA1_DRTYPE) enable((*inhigh*) en115);
        method drvalid(DMA1_DRVALID) enable((*inhigh*) en116);
        method DMA1_RSTN rstn();
    endinterface
    interface Pps7Dma     dma2;
        method aclk(DMA2_ACLK) enable((*inhigh*) en117);
        method daready(DMA2_DAREADY) enable((*inhigh*) en118);
        method DMA2_DATYPE datype();
        method DMA2_DAVALID davalid();
        method drlast(DMA2_DRLAST) enable((*inhigh*) en119);
        method DMA2_DRREADY drready();
        method drtype(DMA2_DRTYPE) enable((*inhigh*) en120);
        method drvalid(DMA2_DRVALID) enable((*inhigh*) en121);
        method DMA2_RSTN rstn();
    endinterface
    interface Pps7Dma     dma3;
        method aclk(DMA3_ACLK) enable((*inhigh*) en122);
        method daready(DMA3_DAREADY) enable((*inhigh*) en123);
        method DMA3_DATYPE datype();
        method DMA3_DAVALID davalid();
        method drlast(DMA3_DRLAST) enable((*inhigh*) en124);
        method DMA3_DRREADY drready();
        method drtype(DMA3_DRTYPE) enable((*inhigh*) en125);
        method drvalid(DMA3_DRVALID) enable((*inhigh*) en126);
        method DMA3_RSTN rstn();
    endinterface
    interface Pps7Enet     enet0;
        method ext_intin(ENET0_EXT_INTIN) enable((*inhigh*) en127);
        method gmii_col(ENET0_GMII_COL) enable((*inhigh*) en128);
        method gmii_crs(ENET0_GMII_CRS) enable((*inhigh*) en129);
        method gmii_rxd(ENET0_GMII_RXD) enable((*inhigh*) en130);
        method gmii_rx_clk(ENET0_GMII_RX_CLK) enable((*inhigh*) en131);
        method gmii_rx_dv(ENET0_GMII_RX_DV) enable((*inhigh*) en132);
        method gmii_rx_er(ENET0_GMII_RX_ER) enable((*inhigh*) en133);
        method ENET0_GMII_TXD gmii_txd();
        method gmii_tx_clk(ENET0_GMII_TX_CLK) enable((*inhigh*) en134);
        method ENET0_GMII_TX_EN gmii_tx_en();
        method ENET0_GMII_TX_ER gmii_tx_er();
        method mdio_i(ENET0_MDIO_I) enable((*inhigh*) en135);
        method ENET0_MDIO_MDC mdio_mdc();
        method ENET0_MDIO_O mdio_o();
        method ENET0_MDIO_T mdio_t();
        method ENET0_PTP_DELAY_REQ_RX ptp_delay_req_rx();
        method ENET0_PTP_DELAY_REQ_TX ptp_delay_req_tx();
        method ENET0_PTP_PDELAY_REQ_RX ptp_pdelay_req_rx();
        method ENET0_PTP_PDELAY_REQ_TX ptp_pdelay_req_tx();
        method ENET0_PTP_PDELAY_RESP_RX ptp_pdelay_resp_rx();
        method ENET0_PTP_PDELAY_RESP_TX ptp_pdelay_resp_tx();
        method ENET0_PTP_SYNC_FRAME_RX ptp_sync_frame_rx();
        method ENET0_PTP_SYNC_FRAME_TX ptp_sync_frame_tx();
        method ENET0_SOF_RX sof_rx();
        method ENET0_SOF_TX sof_tx();
    endinterface
    interface Pps7Enet     enet1;
        method ext_intin(ENET1_EXT_INTIN) enable((*inhigh*) en136);
        method gmii_col(ENET1_GMII_COL) enable((*inhigh*) en137);
        method gmii_crs(ENET1_GMII_CRS) enable((*inhigh*) en138);
        method gmii_rxd(ENET1_GMII_RXD) enable((*inhigh*) en139);
        method gmii_rx_clk(ENET1_GMII_RX_CLK) enable((*inhigh*) en140);
        method gmii_rx_dv(ENET1_GMII_RX_DV) enable((*inhigh*) en141);
        method gmii_rx_er(ENET1_GMII_RX_ER) enable((*inhigh*) en142);
        method ENET1_GMII_TXD gmii_txd();
        method gmii_tx_clk(ENET1_GMII_TX_CLK) enable((*inhigh*) en143);
        method ENET1_GMII_TX_EN gmii_tx_en();
        method ENET1_GMII_TX_ER gmii_tx_er();
        method mdio_i(ENET1_MDIO_I) enable((*inhigh*) en144);
        method ENET1_MDIO_MDC mdio_mdc();
        method ENET1_MDIO_O mdio_o();
        method ENET1_MDIO_T mdio_t();
        method ENET1_PTP_DELAY_REQ_RX ptp_delay_req_rx();
        method ENET1_PTP_DELAY_REQ_TX ptp_delay_req_tx();
        method ENET1_PTP_PDELAY_REQ_RX ptp_pdelay_req_rx();
        method ENET1_PTP_PDELAY_REQ_TX ptp_pdelay_req_tx();
        method ENET1_PTP_PDELAY_RESP_RX ptp_pdelay_resp_rx();
        method ENET1_PTP_PDELAY_RESP_TX ptp_pdelay_resp_tx();
        method ENET1_PTP_SYNC_FRAME_RX ptp_sync_frame_rx();
        method ENET1_PTP_SYNC_FRAME_TX ptp_sync_frame_tx();
        method ENET1_SOF_RX sof_rx();
        method ENET1_SOF_TX sof_tx();
    endinterface
    interface Pps7Event     event_;
        method eventi(EVENT_EVENTI) enable((*inhigh*) en145);
        method EVENT_EVENTO evento();
        method EVENT_STANDBYWFE standbywfe();
        method EVENT_STANDBYWFI standbywfi();
    endinterface
    interface Pps7Fclk     fclk;
        method FCLK_CLK0 clk0();
        method FCLK_CLK1 clk1();
        method FCLK_CLK2 clk2();
        method FCLK_CLK3 clk3();
    endinterface
    interface Pps7Fclk_clktrig     fclk_clktrig0;
        method n(FCLK_CLKTRIG0_N) enable((*inhigh*) en146);
    endinterface
    interface Pps7Fclk_clktrig     fclk_clktrig1;
        method n(FCLK_CLKTRIG1_N) enable((*inhigh*) en147);
    endinterface
    interface Pps7Fclk_clktrig     fclk_clktrig2;
        method n(FCLK_CLKTRIG2_N) enable((*inhigh*) en148);
    endinterface
    interface Pps7Fclk_clktrig     fclk_clktrig3;
        method n(FCLK_CLKTRIG3_N) enable((*inhigh*) en149);
    endinterface
    interface Pps7Fclk_reset     fclk_reset0;
        method FCLK_RESET0_N n();
    endinterface
    interface Pps7Fclk_reset     fclk_reset1;
        method FCLK_RESET1_N n();
    endinterface
    interface Pps7Fclk_reset     fclk_reset2;
        method FCLK_RESET2_N n();
    endinterface
    interface Pps7Fclk_reset     fclk_reset3;
        method FCLK_RESET3_N n();
    endinterface
    interface Pps7Fpga     fpga;
        method idle_n(FPGA_IDLE_N) enable((*inhigh*) en150);
    endinterface
    interface Pps7Ftmd     ftmd;
        method tracein_atid(FTMD_TRACEIN_ATID) enable((*inhigh*) en151);
        method tracein_clk(FTMD_TRACEIN_CLK) enable((*inhigh*) en152);
        method tracein_data(FTMD_TRACEIN_DATA) enable((*inhigh*) en153);
        method tracein_valid(FTMD_TRACEIN_VALID) enable((*inhigh*) en154);
    endinterface
    interface Pps7Ftmt     ftmt;
        method f2p_debug(FTMT_F2P_DEBUG) enable((*inhigh*) en155);
        method f2p_trig(FTMT_F2P_TRIG) enable((*inhigh*) en156);
        method FTMT_F2P_TRIGACK f2p_trigack();
        method FTMT_P2F_DEBUG p2f_debug();
        method FTMT_P2F_TRIG p2f_trig();
        method p2f_trigack(FTMT_P2F_TRIGACK) enable((*inhigh*) en157);
    endinterface
    interface Pps7Gpio     gpio;
        method i(GPIO_I) enable((*inhigh*) en158);
        method GPIO_O o();
        method GPIO_T t();
    endinterface
    interface Pps7I2c     i2c0;
        method scl_i(I2C0_SCL_I) enable((*inhigh*) en159);
        method I2C0_SCL_O scl_o();
        method I2C0_SCL_T scl_t();
        method sda_i(I2C0_SDA_I) enable((*inhigh*) en160);
        method I2C0_SDA_O sda_o();
        method I2C0_SDA_T sda_t();
    endinterface
    interface Pps7I2c     i2c1;
        method scl_i(I2C1_SCL_I) enable((*inhigh*) en161);
        method I2C1_SCL_O scl_o();
        method I2C1_SCL_T scl_t();
        method sda_i(I2C1_SDA_I) enable((*inhigh*) en162);
        method I2C1_SDA_O sda_o();
        method I2C1_SDA_T sda_t();
    endinterface
    interface Pps7Irq     irq;
        method f2p(IRQ_F2P) enable((*inhigh*) en163);
        method IRQ_P2F_CAN0 p2f_can0();
        method IRQ_P2F_CAN1 p2f_can1();
        method IRQ_P2F_CTI p2f_cti();
        method IRQ_P2F_DMAC0 p2f_dmac0();
        method IRQ_P2F_DMAC1 p2f_dmac1();
        method IRQ_P2F_DMAC2 p2f_dmac2();
        method IRQ_P2F_DMAC3 p2f_dmac3();
        method IRQ_P2F_DMAC4 p2f_dmac4();
        method IRQ_P2F_DMAC5 p2f_dmac5();
        method IRQ_P2F_DMAC6 p2f_dmac6();
        method IRQ_P2F_DMAC7 p2f_dmac7();
        method IRQ_P2F_DMAC_ABORT p2f_dmac_abort();
        method IRQ_P2F_ENET0 p2f_enet0();
        method IRQ_P2F_ENET1 p2f_enet1();
        method IRQ_P2F_ENET_WAKE0 p2f_enet_wake0();
        method IRQ_P2F_ENET_WAKE1 p2f_enet_wake1();
        method IRQ_P2F_GPIO p2f_gpio();
        method IRQ_P2F_I2C0 p2f_i2c0();
        method IRQ_P2F_I2C1 p2f_i2c1();
        method IRQ_P2F_QSPI p2f_qspi();
        method IRQ_P2F_SDIO0 p2f_sdio0();
        method IRQ_P2F_SDIO1 p2f_sdio1();
        method IRQ_P2F_SMC p2f_smc();
        method IRQ_P2F_SPI0 p2f_spi0();
        method IRQ_P2F_SPI1 p2f_spi1();
        method IRQ_P2F_UART0 p2f_uart0();
        method IRQ_P2F_UART1 p2f_uart1();
        method IRQ_P2F_USB0 p2f_usb0();
        method IRQ_P2F_USB1 p2f_usb1();
    endinterface
    ifc_inout mio(MIO);
    interface Pps7M_axi_gp     m_axi_gp0;
        method aclk(M_AXI_GP0_ACLK) enable((*inhigh*) en164);
        method M_AXI_GP0_ARADDR araddr();
        method M_AXI_GP0_ARBURST arburst();
        method M_AXI_GP0_ARCACHE arcache();
        method M_AXI_GP0_ARESETN aresetn();
        method M_AXI_GP0_ARID arid();
        method M_AXI_GP0_ARLEN arlen();
        method M_AXI_GP0_ARLOCK arlock();
        method M_AXI_GP0_ARPROT arprot();
        method M_AXI_GP0_ARQOS arqos();
        method arready(M_AXI_GP0_ARREADY) enable((*inhigh*) en165);
        method M_AXI_GP0_ARSIZE arsize();
        method M_AXI_GP0_ARVALID arvalid();
        method M_AXI_GP0_AWADDR awaddr();
        method M_AXI_GP0_AWBURST awburst();
        method M_AXI_GP0_AWCACHE awcache();
        method M_AXI_GP0_AWID awid();
        method M_AXI_GP0_AWLEN awlen();
        method M_AXI_GP0_AWLOCK awlock();
        method M_AXI_GP0_AWPROT awprot();
        method M_AXI_GP0_AWQOS awqos();
        method awready(M_AXI_GP0_AWREADY) enable((*inhigh*) en166);
        method M_AXI_GP0_AWSIZE awsize();
        method M_AXI_GP0_AWVALID awvalid();
        method bid(M_AXI_GP0_BID) enable((*inhigh*) en167);
        method M_AXI_GP0_BREADY bready();
        method bresp(M_AXI_GP0_BRESP) enable((*inhigh*) en168);
        method bvalid(M_AXI_GP0_BVALID) enable((*inhigh*) en169);
        method rdata(M_AXI_GP0_RDATA) enable((*inhigh*) en170);
        method rid(M_AXI_GP0_RID) enable((*inhigh*) en171);
        method rlast(M_AXI_GP0_RLAST) enable((*inhigh*) en172);
        method M_AXI_GP0_RREADY rready();
        method rresp(M_AXI_GP0_RRESP) enable((*inhigh*) en173);
        method rvalid(M_AXI_GP0_RVALID) enable((*inhigh*) en174);
        method M_AXI_GP0_WDATA wdata();
        method M_AXI_GP0_WID wid();
        method M_AXI_GP0_WLAST wlast();
        method wready(M_AXI_GP0_WREADY) enable((*inhigh*) en175);
        method M_AXI_GP0_WSTRB wstrb();
        method M_AXI_GP0_WVALID wvalid();
    endinterface
    interface Pps7M_axi_gp     m_axi_gp1;
        method aclk(M_AXI_GP1_ACLK) enable((*inhigh*) en176);
        method M_AXI_GP1_ARADDR araddr();
        method M_AXI_GP1_ARBURST arburst();
        method M_AXI_GP1_ARCACHE arcache();
        method M_AXI_GP1_ARESETN aresetn();
        method M_AXI_GP1_ARID arid();
        method M_AXI_GP1_ARLEN arlen();
        method M_AXI_GP1_ARLOCK arlock();
        method M_AXI_GP1_ARPROT arprot();
        method M_AXI_GP1_ARQOS arqos();
        method arready(M_AXI_GP1_ARREADY) enable((*inhigh*) en177);
        method M_AXI_GP1_ARSIZE arsize();
        method M_AXI_GP1_ARVALID arvalid();
        method M_AXI_GP1_AWADDR awaddr();
        method M_AXI_GP1_AWBURST awburst();
        method M_AXI_GP1_AWCACHE awcache();
        method M_AXI_GP1_AWID awid();
        method M_AXI_GP1_AWLEN awlen();
        method M_AXI_GP1_AWLOCK awlock();
        method M_AXI_GP1_AWPROT awprot();
        method M_AXI_GP1_AWQOS awqos();
        method awready(M_AXI_GP1_AWREADY) enable((*inhigh*) en178);
        method M_AXI_GP1_AWSIZE awsize();
        method M_AXI_GP1_AWVALID awvalid();
        method bid(M_AXI_GP1_BID) enable((*inhigh*) en179);
        method M_AXI_GP1_BREADY bready();
        method bresp(M_AXI_GP1_BRESP) enable((*inhigh*) en180);
        method bvalid(M_AXI_GP1_BVALID) enable((*inhigh*) en181);
        method rdata(M_AXI_GP1_RDATA) enable((*inhigh*) en182);
        method rid(M_AXI_GP1_RID) enable((*inhigh*) en183);
        method rlast(M_AXI_GP1_RLAST) enable((*inhigh*) en184);
        method M_AXI_GP1_RREADY rready();
        method rresp(M_AXI_GP1_RRESP) enable((*inhigh*) en185);
        method rvalid(M_AXI_GP1_RVALID) enable((*inhigh*) en186);
        method M_AXI_GP1_WDATA wdata();
        method M_AXI_GP1_WID wid();
        method M_AXI_GP1_WLAST wlast();
        method wready(M_AXI_GP1_WREADY) enable((*inhigh*) en187);
        method M_AXI_GP1_WSTRB wstrb();
        method M_AXI_GP1_WVALID wvalid();
    endinterface
    interface Pps7Pjtag     pjtag;
        method tck(PJTAG_TCK) enable((*inhigh*) en188);
        method td_i(PJTAG_TD_I) enable((*inhigh*) en189);
        method PJTAG_TD_O td_o();
        method PJTAG_TD_T td_t();
        method tms(PJTAG_TMS) enable((*inhigh*) en190);
    endinterface
    interface Pps7Ps     ps;
        method clk(PS_CLK) enable((*inhigh*) en191);
        method porb(PS_PORB) enable((*inhigh*) en192);
        method srstb(PS_SRSTB) enable((*inhigh*) en193);
    endinterface
    interface Pps7Sdio     sdio0;
        method SDIO0_BUSPOW buspow();
        method SDIO0_BUSVOLT busvolt();
        method cdn(SDIO0_CDN) enable((*inhigh*) en194);
        method SDIO0_CLK clk();
        method clk_fb(SDIO0_CLK_FB) enable((*inhigh*) en195);
        method cmd_i(SDIO0_CMD_I) enable((*inhigh*) en196);
        method SDIO0_CMD_O cmd_o();
        method SDIO0_CMD_T cmd_t();
        method data_i(SDIO0_DATA_I) enable((*inhigh*) en197);
        method SDIO0_DATA_O data_o();
        method SDIO0_DATA_T data_t();
        method SDIO0_LED led();
        method wp(SDIO0_WP) enable((*inhigh*) en198);
    endinterface
    interface Pps7Sdio     sdio1;
        method SDIO1_BUSPOW buspow();
        method SDIO1_BUSVOLT busvolt();
        method cdn(SDIO1_CDN) enable((*inhigh*) en199);
        method SDIO1_CLK clk();
        method clk_fb(SDIO1_CLK_FB) enable((*inhigh*) en200);
        method cmd_i(SDIO1_CMD_I) enable((*inhigh*) en201);
        method SDIO1_CMD_O cmd_o();
        method SDIO1_CMD_T cmd_t();
        method data_i(SDIO1_DATA_I) enable((*inhigh*) en202);
        method SDIO1_DATA_O data_o();
        method SDIO1_DATA_T data_t();
        method SDIO1_LED led();
        method wp(SDIO1_WP) enable((*inhigh*) en203);
    endinterface
    interface Pps7Spi     spi0;
        method miso_i(SPI0_MISO_I) enable((*inhigh*) en204);
        method SPI0_MISO_O miso_o();
        method SPI0_MISO_T miso_t();
        method mosi_i(SPI0_MOSI_I) enable((*inhigh*) en205);
        method SPI0_MOSI_O mosi_o();
        method SPI0_MOSI_T mosi_t();
        method sclk_i(SPI0_SCLK_I) enable((*inhigh*) en206);
        method SPI0_SCLK_O sclk_o();
        method SPI0_SCLK_T sclk_t();
        method SPI0_SS1_O ss1_o();
        method SPI0_SS2_O ss2_o();
        method ss_i(SPI0_SS_I) enable((*inhigh*) en207);
        method SPI0_SS_O ss_o();
        method SPI0_SS_T ss_t();
    endinterface
    interface Pps7Spi     spi1;
        method miso_i(SPI1_MISO_I) enable((*inhigh*) en208);
        method SPI1_MISO_O miso_o();
        method SPI1_MISO_T miso_t();
        method mosi_i(SPI1_MOSI_I) enable((*inhigh*) en209);
        method SPI1_MOSI_O mosi_o();
        method SPI1_MOSI_T mosi_t();
        method sclk_i(SPI1_SCLK_I) enable((*inhigh*) en210);
        method SPI1_SCLK_O sclk_o();
        method SPI1_SCLK_T sclk_t();
        method SPI1_SS1_O ss1_o();
        method SPI1_SS2_O ss2_o();
        method ss_i(SPI1_SS_I) enable((*inhigh*) en211);
        method SPI1_SS_O ss_o();
        method SPI1_SS_T ss_t();
    endinterface
    interface Pps7Sram     sram;
        method intin(SRAM_INTIN) enable((*inhigh*) en212);
    endinterface
    interface Pps7S_axi_acp     s_axi_acp;
        method aclk(S_AXI_ACP_ACLK) enable((*inhigh*) en213);
        method araddr(S_AXI_ACP_ARADDR) enable((*inhigh*) en214);
        method arburst(S_AXI_ACP_ARBURST) enable((*inhigh*) en215);
        method arcache(S_AXI_ACP_ARCACHE) enable((*inhigh*) en216);
        method S_AXI_ACP_ARESETN aresetn();
        method arid(S_AXI_ACP_ARID) enable((*inhigh*) en217);
        method arlen(S_AXI_ACP_ARLEN) enable((*inhigh*) en218);
        method arlock(S_AXI_ACP_ARLOCK) enable((*inhigh*) en219);
        method arprot(S_AXI_ACP_ARPROT) enable((*inhigh*) en220);
        method arqos(S_AXI_ACP_ARQOS) enable((*inhigh*) en221);
        method S_AXI_ACP_ARREADY arready();
        method arsize(S_AXI_ACP_ARSIZE) enable((*inhigh*) en222);
        method aruser(S_AXI_ACP_ARUSER) enable((*inhigh*) en223);
        method arvalid(S_AXI_ACP_ARVALID) enable((*inhigh*) en224);
        method awaddr(S_AXI_ACP_AWADDR) enable((*inhigh*) en225);
        method awburst(S_AXI_ACP_AWBURST) enable((*inhigh*) en226);
        method awcache(S_AXI_ACP_AWCACHE) enable((*inhigh*) en227);
        method awid(S_AXI_ACP_AWID) enable((*inhigh*) en228);
        method awlen(S_AXI_ACP_AWLEN) enable((*inhigh*) en229);
        method awlock(S_AXI_ACP_AWLOCK) enable((*inhigh*) en230);
        method awprot(S_AXI_ACP_AWPROT) enable((*inhigh*) en231);
        method awqos(S_AXI_ACP_AWQOS) enable((*inhigh*) en232);
        method S_AXI_ACP_AWREADY awready();
        method awsize(S_AXI_ACP_AWSIZE) enable((*inhigh*) en233);
        method awuser(S_AXI_ACP_AWUSER) enable((*inhigh*) en234);
        method awvalid(S_AXI_ACP_AWVALID) enable((*inhigh*) en235);
        method S_AXI_ACP_BID bid();
        method bready(S_AXI_ACP_BREADY) enable((*inhigh*) en236);
        method S_AXI_ACP_BRESP bresp();
        method S_AXI_ACP_BVALID bvalid();
        method S_AXI_ACP_RDATA rdata();
        method S_AXI_ACP_RID rid();
        method S_AXI_ACP_RLAST rlast();
        method rready(S_AXI_ACP_RREADY) enable((*inhigh*) en237);
        method S_AXI_ACP_RRESP rresp();
        method S_AXI_ACP_RVALID rvalid();
        method wdata(S_AXI_ACP_WDATA) enable((*inhigh*) en238);
        method wid(S_AXI_ACP_WID) enable((*inhigh*) en239);
        method wlast(S_AXI_ACP_WLAST) enable((*inhigh*) en240);
        method S_AXI_ACP_WREADY wready();
        method wstrb(S_AXI_ACP_WSTRB) enable((*inhigh*) en241);
        method wvalid(S_AXI_ACP_WVALID) enable((*inhigh*) en242);
    endinterface
    interface Pps7S_axi_gp     s_axi_gp0;
        method aclk(S_AXI_GP0_ACLK) enable((*inhigh*) en243);
        method araddr(S_AXI_GP0_ARADDR) enable((*inhigh*) en244);
        method arburst(S_AXI_GP0_ARBURST) enable((*inhigh*) en245);
        method arcache(S_AXI_GP0_ARCACHE) enable((*inhigh*) en246);
        method S_AXI_GP0_ARESETN aresetn();
        method arid(S_AXI_GP0_ARID) enable((*inhigh*) en247);
        method arlen(S_AXI_GP0_ARLEN) enable((*inhigh*) en248);
        method arlock(S_AXI_GP0_ARLOCK) enable((*inhigh*) en249);
        method arprot(S_AXI_GP0_ARPROT) enable((*inhigh*) en250);
        method arqos(S_AXI_GP0_ARQOS) enable((*inhigh*) en251);
        method S_AXI_GP0_ARREADY arready();
        method arsize(S_AXI_GP0_ARSIZE) enable((*inhigh*) en252);
        method arvalid(S_AXI_GP0_ARVALID) enable((*inhigh*) en253);
        method awaddr(S_AXI_GP0_AWADDR) enable((*inhigh*) en254);
        method awburst(S_AXI_GP0_AWBURST) enable((*inhigh*) en255);
        method awcache(S_AXI_GP0_AWCACHE) enable((*inhigh*) en256);
        method awid(S_AXI_GP0_AWID) enable((*inhigh*) en257);
        method awlen(S_AXI_GP0_AWLEN) enable((*inhigh*) en258);
        method awlock(S_AXI_GP0_AWLOCK) enable((*inhigh*) en259);
        method awprot(S_AXI_GP0_AWPROT) enable((*inhigh*) en260);
        method awqos(S_AXI_GP0_AWQOS) enable((*inhigh*) en261);
        method S_AXI_GP0_AWREADY awready();
        method awsize(S_AXI_GP0_AWSIZE) enable((*inhigh*) en262);
        method awvalid(S_AXI_GP0_AWVALID) enable((*inhigh*) en263);
        method S_AXI_GP0_BID bid();
        method bready(S_AXI_GP0_BREADY) enable((*inhigh*) en264);
        method S_AXI_GP0_BRESP bresp();
        method S_AXI_GP0_BVALID bvalid();
        method S_AXI_GP0_RDATA rdata();
        method S_AXI_GP0_RID rid();
        method S_AXI_GP0_RLAST rlast();
        method rready(S_AXI_GP0_RREADY) enable((*inhigh*) en265);
        method S_AXI_GP0_RRESP rresp();
        method S_AXI_GP0_RVALID rvalid();
        method wdata(S_AXI_GP0_WDATA) enable((*inhigh*) en266);
        method wid(S_AXI_GP0_WID) enable((*inhigh*) en267);
        method wlast(S_AXI_GP0_WLAST) enable((*inhigh*) en268);
        method S_AXI_GP0_WREADY wready();
        method wstrb(S_AXI_GP0_WSTRB) enable((*inhigh*) en269);
        method wvalid(S_AXI_GP0_WVALID) enable((*inhigh*) en270);
    endinterface
    interface Pps7S_axi_gp     s_axi_gp1;
        method aclk(S_AXI_GP1_ACLK) enable((*inhigh*) en271);
        method araddr(S_AXI_GP1_ARADDR) enable((*inhigh*) en272);
        method arburst(S_AXI_GP1_ARBURST) enable((*inhigh*) en273);
        method arcache(S_AXI_GP1_ARCACHE) enable((*inhigh*) en274);
        method S_AXI_GP1_ARESETN aresetn();
        method arid(S_AXI_GP1_ARID) enable((*inhigh*) en275);
        method arlen(S_AXI_GP1_ARLEN) enable((*inhigh*) en276);
        method arlock(S_AXI_GP1_ARLOCK) enable((*inhigh*) en277);
        method arprot(S_AXI_GP1_ARPROT) enable((*inhigh*) en278);
        method arqos(S_AXI_GP1_ARQOS) enable((*inhigh*) en279);
        method S_AXI_GP1_ARREADY arready();
        method arsize(S_AXI_GP1_ARSIZE) enable((*inhigh*) en280);
        method arvalid(S_AXI_GP1_ARVALID) enable((*inhigh*) en281);
        method awaddr(S_AXI_GP1_AWADDR) enable((*inhigh*) en282);
        method awburst(S_AXI_GP1_AWBURST) enable((*inhigh*) en283);
        method awcache(S_AXI_GP1_AWCACHE) enable((*inhigh*) en284);
        method awid(S_AXI_GP1_AWID) enable((*inhigh*) en285);
        method awlen(S_AXI_GP1_AWLEN) enable((*inhigh*) en286);
        method awlock(S_AXI_GP1_AWLOCK) enable((*inhigh*) en287);
        method awprot(S_AXI_GP1_AWPROT) enable((*inhigh*) en288);
        method awqos(S_AXI_GP1_AWQOS) enable((*inhigh*) en289);
        method S_AXI_GP1_AWREADY awready();
        method awsize(S_AXI_GP1_AWSIZE) enable((*inhigh*) en290);
        method awvalid(S_AXI_GP1_AWVALID) enable((*inhigh*) en291);
        method S_AXI_GP1_BID bid();
        method bready(S_AXI_GP1_BREADY) enable((*inhigh*) en292);
        method S_AXI_GP1_BRESP bresp();
        method S_AXI_GP1_BVALID bvalid();
        method S_AXI_GP1_RDATA rdata();
        method S_AXI_GP1_RID rid();
        method S_AXI_GP1_RLAST rlast();
        method rready(S_AXI_GP1_RREADY) enable((*inhigh*) en293);
        method S_AXI_GP1_RRESP rresp();
        method S_AXI_GP1_RVALID rvalid();
        method wdata(S_AXI_GP1_WDATA) enable((*inhigh*) en294);
        method wid(S_AXI_GP1_WID) enable((*inhigh*) en295);
        method wlast(S_AXI_GP1_WLAST) enable((*inhigh*) en296);
        method S_AXI_GP1_WREADY wready();
        method wstrb(S_AXI_GP1_WSTRB) enable((*inhigh*) en297);
        method wvalid(S_AXI_GP1_WVALID) enable((*inhigh*) en298);
    endinterface
    interface Pps7S_axi_hp     s_axi_hp0;
        method aclk(S_AXI_HP0_ACLK) enable((*inhigh*) en299);
        method araddr(S_AXI_HP0_ARADDR) enable((*inhigh*) en300);
        method arburst(S_AXI_HP0_ARBURST) enable((*inhigh*) en301);
        method arcache(S_AXI_HP0_ARCACHE) enable((*inhigh*) en302);
        method S_AXI_HP0_ARESETN aresetn();
        method arid(S_AXI_HP0_ARID) enable((*inhigh*) en303);
        method arlen(S_AXI_HP0_ARLEN) enable((*inhigh*) en304);
        method arlock(S_AXI_HP0_ARLOCK) enable((*inhigh*) en305);
        method arprot(S_AXI_HP0_ARPROT) enable((*inhigh*) en306);
        method arqos(S_AXI_HP0_ARQOS) enable((*inhigh*) en307);
        method S_AXI_HP0_ARREADY arready();
        method arsize(S_AXI_HP0_ARSIZE) enable((*inhigh*) en308);
        method arvalid(S_AXI_HP0_ARVALID) enable((*inhigh*) en309);
        method awaddr(S_AXI_HP0_AWADDR) enable((*inhigh*) en310);
        method awburst(S_AXI_HP0_AWBURST) enable((*inhigh*) en311);
        method awcache(S_AXI_HP0_AWCACHE) enable((*inhigh*) en312);
        method awid(S_AXI_HP0_AWID) enable((*inhigh*) en313);
        method awlen(S_AXI_HP0_AWLEN) enable((*inhigh*) en314);
        method awlock(S_AXI_HP0_AWLOCK) enable((*inhigh*) en315);
        method awprot(S_AXI_HP0_AWPROT) enable((*inhigh*) en316);
        method awqos(S_AXI_HP0_AWQOS) enable((*inhigh*) en317);
        method S_AXI_HP0_AWREADY awready();
        method awsize(S_AXI_HP0_AWSIZE) enable((*inhigh*) en318);
        method awvalid(S_AXI_HP0_AWVALID) enable((*inhigh*) en319);
        method S_AXI_HP0_BID bid();
        method bready(S_AXI_HP0_BREADY) enable((*inhigh*) en320);
        method S_AXI_HP0_BRESP bresp();
        method S_AXI_HP0_BVALID bvalid();
        method S_AXI_HP0_RACOUNT racount();
        method S_AXI_HP0_RCOUNT rcount();
        method S_AXI_HP0_RDATA rdata();
        method rdissuecap1_en(S_AXI_HP0_RDISSUECAP1_EN) enable((*inhigh*) en321);
        method S_AXI_HP0_RID rid();
        method S_AXI_HP0_RLAST rlast();
        method rready(S_AXI_HP0_RREADY) enable((*inhigh*) en322);
        method S_AXI_HP0_RRESP rresp();
        method S_AXI_HP0_RVALID rvalid();
        method S_AXI_HP0_WACOUNT wacount();
        method S_AXI_HP0_WCOUNT wcount();
        method wdata(S_AXI_HP0_WDATA) enable((*inhigh*) en323);
        method wid(S_AXI_HP0_WID) enable((*inhigh*) en324);
        method wlast(S_AXI_HP0_WLAST) enable((*inhigh*) en325);
        method S_AXI_HP0_WREADY wready();
        method wrissuecap1_en(S_AXI_HP0_WRISSUECAP1_EN) enable((*inhigh*) en326);
        method wstrb(S_AXI_HP0_WSTRB) enable((*inhigh*) en327);
        method wvalid(S_AXI_HP0_WVALID) enable((*inhigh*) en328);
    endinterface
    interface Pps7S_axi_hp     s_axi_hp1;
        method aclk(S_AXI_HP1_ACLK) enable((*inhigh*) en329);
        method araddr(S_AXI_HP1_ARADDR) enable((*inhigh*) en330);
        method arburst(S_AXI_HP1_ARBURST) enable((*inhigh*) en331);
        method arcache(S_AXI_HP1_ARCACHE) enable((*inhigh*) en332);
        method S_AXI_HP1_ARESETN aresetn();
        method arid(S_AXI_HP1_ARID) enable((*inhigh*) en333);
        method arlen(S_AXI_HP1_ARLEN) enable((*inhigh*) en334);
        method arlock(S_AXI_HP1_ARLOCK) enable((*inhigh*) en335);
        method arprot(S_AXI_HP1_ARPROT) enable((*inhigh*) en336);
        method arqos(S_AXI_HP1_ARQOS) enable((*inhigh*) en337);
        method S_AXI_HP1_ARREADY arready();
        method arsize(S_AXI_HP1_ARSIZE) enable((*inhigh*) en338);
        method arvalid(S_AXI_HP1_ARVALID) enable((*inhigh*) en339);
        method awaddr(S_AXI_HP1_AWADDR) enable((*inhigh*) en340);
        method awburst(S_AXI_HP1_AWBURST) enable((*inhigh*) en341);
        method awcache(S_AXI_HP1_AWCACHE) enable((*inhigh*) en342);
        method awid(S_AXI_HP1_AWID) enable((*inhigh*) en343);
        method awlen(S_AXI_HP1_AWLEN) enable((*inhigh*) en344);
        method awlock(S_AXI_HP1_AWLOCK) enable((*inhigh*) en345);
        method awprot(S_AXI_HP1_AWPROT) enable((*inhigh*) en346);
        method awqos(S_AXI_HP1_AWQOS) enable((*inhigh*) en347);
        method S_AXI_HP1_AWREADY awready();
        method awsize(S_AXI_HP1_AWSIZE) enable((*inhigh*) en348);
        method awvalid(S_AXI_HP1_AWVALID) enable((*inhigh*) en349);
        method S_AXI_HP1_BID bid();
        method bready(S_AXI_HP1_BREADY) enable((*inhigh*) en350);
        method S_AXI_HP1_BRESP bresp();
        method S_AXI_HP1_BVALID bvalid();
        method S_AXI_HP1_RACOUNT racount();
        method S_AXI_HP1_RCOUNT rcount();
        method S_AXI_HP1_RDATA rdata();
        method rdissuecap1_en(S_AXI_HP1_RDISSUECAP1_EN) enable((*inhigh*) en351);
        method S_AXI_HP1_RID rid();
        method S_AXI_HP1_RLAST rlast();
        method rready(S_AXI_HP1_RREADY) enable((*inhigh*) en352);
        method S_AXI_HP1_RRESP rresp();
        method S_AXI_HP1_RVALID rvalid();
        method S_AXI_HP1_WACOUNT wacount();
        method S_AXI_HP1_WCOUNT wcount();
        method wdata(S_AXI_HP1_WDATA) enable((*inhigh*) en353);
        method wid(S_AXI_HP1_WID) enable((*inhigh*) en354);
        method wlast(S_AXI_HP1_WLAST) enable((*inhigh*) en355);
        method S_AXI_HP1_WREADY wready();
        method wrissuecap1_en(S_AXI_HP1_WRISSUECAP1_EN) enable((*inhigh*) en356);
        method wstrb(S_AXI_HP1_WSTRB) enable((*inhigh*) en357);
        method wvalid(S_AXI_HP1_WVALID) enable((*inhigh*) en358);
    endinterface
    interface Pps7S_axi_hp     s_axi_hp2;
        method aclk(S_AXI_HP2_ACLK) enable((*inhigh*) en359);
        method araddr(S_AXI_HP2_ARADDR) enable((*inhigh*) en360);
        method arburst(S_AXI_HP2_ARBURST) enable((*inhigh*) en361);
        method arcache(S_AXI_HP2_ARCACHE) enable((*inhigh*) en362);
        method S_AXI_HP2_ARESETN aresetn();
        method arid(S_AXI_HP2_ARID) enable((*inhigh*) en363);
        method arlen(S_AXI_HP2_ARLEN) enable((*inhigh*) en364);
        method arlock(S_AXI_HP2_ARLOCK) enable((*inhigh*) en365);
        method arprot(S_AXI_HP2_ARPROT) enable((*inhigh*) en366);
        method arqos(S_AXI_HP2_ARQOS) enable((*inhigh*) en367);
        method S_AXI_HP2_ARREADY arready();
        method arsize(S_AXI_HP2_ARSIZE) enable((*inhigh*) en368);
        method arvalid(S_AXI_HP2_ARVALID) enable((*inhigh*) en369);
        method awaddr(S_AXI_HP2_AWADDR) enable((*inhigh*) en370);
        method awburst(S_AXI_HP2_AWBURST) enable((*inhigh*) en371);
        method awcache(S_AXI_HP2_AWCACHE) enable((*inhigh*) en372);
        method awid(S_AXI_HP2_AWID) enable((*inhigh*) en373);
        method awlen(S_AXI_HP2_AWLEN) enable((*inhigh*) en374);
        method awlock(S_AXI_HP2_AWLOCK) enable((*inhigh*) en375);
        method awprot(S_AXI_HP2_AWPROT) enable((*inhigh*) en376);
        method awqos(S_AXI_HP2_AWQOS) enable((*inhigh*) en377);
        method S_AXI_HP2_AWREADY awready();
        method awsize(S_AXI_HP2_AWSIZE) enable((*inhigh*) en378);
        method awvalid(S_AXI_HP2_AWVALID) enable((*inhigh*) en379);
        method S_AXI_HP2_BID bid();
        method bready(S_AXI_HP2_BREADY) enable((*inhigh*) en380);
        method S_AXI_HP2_BRESP bresp();
        method S_AXI_HP2_BVALID bvalid();
        method S_AXI_HP2_RACOUNT racount();
        method S_AXI_HP2_RCOUNT rcount();
        method S_AXI_HP2_RDATA rdata();
        method rdissuecap1_en(S_AXI_HP2_RDISSUECAP1_EN) enable((*inhigh*) en381);
        method S_AXI_HP2_RID rid();
        method S_AXI_HP2_RLAST rlast();
        method rready(S_AXI_HP2_RREADY) enable((*inhigh*) en382);
        method S_AXI_HP2_RRESP rresp();
        method S_AXI_HP2_RVALID rvalid();
        method S_AXI_HP2_WACOUNT wacount();
        method S_AXI_HP2_WCOUNT wcount();
        method wdata(S_AXI_HP2_WDATA) enable((*inhigh*) en383);
        method wid(S_AXI_HP2_WID) enable((*inhigh*) en384);
        method wlast(S_AXI_HP2_WLAST) enable((*inhigh*) en385);
        method S_AXI_HP2_WREADY wready();
        method wrissuecap1_en(S_AXI_HP2_WRISSUECAP1_EN) enable((*inhigh*) en386);
        method wstrb(S_AXI_HP2_WSTRB) enable((*inhigh*) en387);
        method wvalid(S_AXI_HP2_WVALID) enable((*inhigh*) en388);
    endinterface
    interface Pps7S_axi_hp     s_axi_hp3;
        method aclk(S_AXI_HP3_ACLK) enable((*inhigh*) en389);
        method araddr(S_AXI_HP3_ARADDR) enable((*inhigh*) en390);
        method arburst(S_AXI_HP3_ARBURST) enable((*inhigh*) en391);
        method arcache(S_AXI_HP3_ARCACHE) enable((*inhigh*) en392);
        method S_AXI_HP3_ARESETN aresetn();
        method arid(S_AXI_HP3_ARID) enable((*inhigh*) en393);
        method arlen(S_AXI_HP3_ARLEN) enable((*inhigh*) en394);
        method arlock(S_AXI_HP3_ARLOCK) enable((*inhigh*) en395);
        method arprot(S_AXI_HP3_ARPROT) enable((*inhigh*) en396);
        method arqos(S_AXI_HP3_ARQOS) enable((*inhigh*) en397);
        method S_AXI_HP3_ARREADY arready();
        method arsize(S_AXI_HP3_ARSIZE) enable((*inhigh*) en398);
        method arvalid(S_AXI_HP3_ARVALID) enable((*inhigh*) en399);
        method awaddr(S_AXI_HP3_AWADDR) enable((*inhigh*) en400);
        method awburst(S_AXI_HP3_AWBURST) enable((*inhigh*) en401);
        method awcache(S_AXI_HP3_AWCACHE) enable((*inhigh*) en402);
        method awid(S_AXI_HP3_AWID) enable((*inhigh*) en403);
        method awlen(S_AXI_HP3_AWLEN) enable((*inhigh*) en404);
        method awlock(S_AXI_HP3_AWLOCK) enable((*inhigh*) en405);
        method awprot(S_AXI_HP3_AWPROT) enable((*inhigh*) en406);
        method awqos(S_AXI_HP3_AWQOS) enable((*inhigh*) en407);
        method S_AXI_HP3_AWREADY awready();
        method awsize(S_AXI_HP3_AWSIZE) enable((*inhigh*) en408);
        method awvalid(S_AXI_HP3_AWVALID) enable((*inhigh*) en409);
        method S_AXI_HP3_BID bid();
        method bready(S_AXI_HP3_BREADY) enable((*inhigh*) en410);
        method S_AXI_HP3_BRESP bresp();
        method S_AXI_HP3_BVALID bvalid();
        method S_AXI_HP3_RACOUNT racount();
        method S_AXI_HP3_RCOUNT rcount();
        method S_AXI_HP3_RDATA rdata();
        method rdissuecap1_en(S_AXI_HP3_RDISSUECAP1_EN) enable((*inhigh*) en411);
        method S_AXI_HP3_RID rid();
        method S_AXI_HP3_RLAST rlast();
        method rready(S_AXI_HP3_RREADY) enable((*inhigh*) en412);
        method S_AXI_HP3_RRESP rresp();
        method S_AXI_HP3_RVALID rvalid();
        method S_AXI_HP3_WACOUNT wacount();
        method S_AXI_HP3_WCOUNT wcount();
        method wdata(S_AXI_HP3_WDATA) enable((*inhigh*) en413);
        method wid(S_AXI_HP3_WID) enable((*inhigh*) en414);
        method wlast(S_AXI_HP3_WLAST) enable((*inhigh*) en415);
        method S_AXI_HP3_WREADY wready();
        method wrissuecap1_en(S_AXI_HP3_WRISSUECAP1_EN) enable((*inhigh*) en416);
        method wstrb(S_AXI_HP3_WSTRB) enable((*inhigh*) en417);
        method wvalid(S_AXI_HP3_WVALID) enable((*inhigh*) en418);
    endinterface
    interface Pps7Trace     trace;
        method clk(TRACE_CLK) enable((*inhigh*) en419);
        method TRACE_CTL ctl();
        method TRACE_DATA data();
    endinterface
    interface Pps7Ttc     ttc0;
        method clk0_in(TTC0_CLK0_IN) enable((*inhigh*) en420);
        method clk1_in(TTC0_CLK1_IN) enable((*inhigh*) en421);
        method clk2_in(TTC0_CLK2_IN) enable((*inhigh*) en422);
        method TTC0_WAVE0_OUT wave0_out();
        method TTC0_WAVE1_OUT wave1_out();
        method TTC0_WAVE2_OUT wave2_out();
    endinterface
    interface Pps7Ttc     ttc1;
        method clk0_in(TTC1_CLK0_IN) enable((*inhigh*) en423);
        method clk1_in(TTC1_CLK1_IN) enable((*inhigh*) en424);
        method clk2_in(TTC1_CLK2_IN) enable((*inhigh*) en425);
        method TTC1_WAVE0_OUT wave0_out();
        method TTC1_WAVE1_OUT wave1_out();
        method TTC1_WAVE2_OUT wave2_out();
    endinterface
    interface Pps7Uart     uart0;
        method ctsn(UART0_CTSN) enable((*inhigh*) en426);
        method dcdn(UART0_DCDN) enable((*inhigh*) en427);
        method dsrn(UART0_DSRN) enable((*inhigh*) en428);
        method UART0_DTRN dtrn();
        method rin(UART0_RIN) enable((*inhigh*) en429);
        method UART0_RTSN rtsn();
        method rx(UART0_RX) enable((*inhigh*) en430);
        method UART0_TX tx();
    endinterface
    interface Pps7Uart     uart1;
        method ctsn(UART1_CTSN) enable((*inhigh*) en431);
        method dcdn(UART1_DCDN) enable((*inhigh*) en432);
        method dsrn(UART1_DSRN) enable((*inhigh*) en433);
        method UART1_DTRN dtrn();
        method rin(UART1_RIN) enable((*inhigh*) en434);
        method UART1_RTSN rtsn();
        method rx(UART1_RX) enable((*inhigh*) en435);
        method UART1_TX tx();
    endinterface
    interface Pps7Usb     usb0;
        method USB0_PORT_INDCTL port_indctl();
        method vbus_pwrfault(USB0_VBUS_PWRFAULT) enable((*inhigh*) en436);
        method USB0_VBUS_PWRSELECT vbus_pwrselect();
    endinterface
    interface Pps7Usb     usb1;
        method USB1_PORT_INDCTL port_indctl();
        method vbus_pwrfault(USB1_VBUS_PWRFAULT) enable((*inhigh*) en437);
        method USB1_VBUS_PWRSELECT vbus_pwrselect();
    endinterface
    interface Pps7Wdt     wdt;
        method clk_in(WDT_CLK_IN) enable((*inhigh*) en438);
        method WDT_RST_OUT rst_out();
    endinterface
endmodule
