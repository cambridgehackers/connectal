// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;
import BRAM::*;
import DefaultValue::*;
import Connectable::*;

// portz libraries
import Leds::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import PortalMemory::*;
import MemTypes::*;
import MemServer::*;
import MemServerInternal::*;
import SGList::*;


// generated by tool
import NandSimRequestWrapper::*;
import DmaDebugRequestWrapper::*;
import SGListConfigRequestWrapper::*;
import StrstrRequestWrapper::*;

import NandSimIndicationProxy::*;
import DmaDebugIndicationProxy::*;
import SGListConfigIndicationProxy::*;
import StrstrIndicationProxy::*;

// defined by user
import NandSim::*;
import NandSimNames::*;
import Strstr::*;

module mkPortalTop(StdPortalDmaTop#(PhysAddrWidth));
   
   // nandsim 
   NandSimIndicationProxy nandSimIndicationProxy <- mkNandSimIndicationProxy(NandSimIndication);
   NandSim nandSim <- mkNandSim(nandSimIndicationProxy.ifc);
   NandSimRequestWrapper nandSimRequestWrapper <- mkNandSimRequestWrapper(NandSimRequest,nandSim.request);
   
   // strstr algo
   StrstrIndicationProxy strstrIndicationProxy <- mkStrstrIndicationProxy(AlgoIndication);
   Strstr#(1,64) strstr <- mkStrstr(strstrIndicationProxy.ifc);
   StrstrRequestWrapper strstrRequestWrapper <- mkStrstrRequestWrapper(AlgoRequest,strstr.request);
   
   // backing store sglist
   SGListConfigIndicationProxy backingStoreSGListConfigIndicationProxy <- mkSGListConfigIndicationProxy(BackingStoreSGListConfigIndication);
   SGListMMU#(PhysAddrWidth) backingStoreSGList <- mkSGListMMU(0, True, backingStoreSGListConfigIndicationProxy.ifc);
   SGListConfigRequestWrapper backingStoreSGListConfigRequestWrapper <- mkSGListConfigRequestWrapper(BackingStoreSGListConfigRequest, backingStoreSGList.request);

   // algo sglist
   SGListConfigIndicationProxy algoSGListConfigIndicationProxy <- mkSGListConfigIndicationProxy(AlgoSGListConfigIndication);
   SGListMMU#(PhysAddrWidth) algoSGList <- mkSGListMMU(1, True, algoSGListConfigIndicationProxy.ifc);
   SGListConfigRequestWrapper algoSGListConfigRequestWrapper <- mkSGListConfigRequestWrapper(AlgoSGListConfigRequest, algoSGList.request);
   
   // nandsim sglist
   SGListConfigIndicationProxy nandsimSGListConfigIndicationProxy <- mkSGListConfigIndicationProxy(NandsimSGListConfigIndication);
   SGListMMU#(PhysAddrWidth) nandsimSGList <- mkSGListMMU(0, False, nandsimSGListConfigIndicationProxy.ifc);
   SGListConfigRequestWrapper nandsimSGListConfigRequestWrapper <- mkSGListConfigRequestWrapper(NandsimSGListConfigRequest, nandsimSGList.request);
   
   // host memory dma server
   DmaDebugIndicationProxy hostDmaDebugIndicationProxy <- mkDmaDebugIndicationProxy(HostmemDmaDebugIndication);
   let rcs = cons(strstr.config_read_client,cons(nandSim.readClient, nil));
   MemServer#(PhysAddrWidth,64,1) hostDma <- mkMemServerRW(hostDmaDebugIndicationProxy.ifc, rcs, cons(nandSim.writeClient, nil), cons(backingStoreSGList,cons(algoSGList,nil)));
   DmaDebugRequestWrapper hostDmaDebugRequestWrapper <- mkDmaDebugRequestWrapper(HostmemDmaDebugRequest, hostDma.request);

   // nandsim memory dma server
   DmaDebugIndicationProxy nandsimDmaDebugIndicationProxy <- mkDmaDebugIndicationProxy(NandsimDmaDebugIndication);   
   MemServer#(PhysAddrWidth,64,1) nandsimDma <- mkMemServerR(nandsimDmaDebugIndicationProxy.ifc, cons(strstr.haystack_read_client,nil), cons(nandsimSGList,nil));
   DmaDebugRequestWrapper nandsimDmaRequestWrapper <- mkDmaDebugRequestWrapper(NandsimDmaDebugRequest, nandsimDma.request);
   mkConnection(nandsimDma.masters[0], nandSim.memSlave);
   
   Vector#(14,StdPortal) portals;

   portals[0] = nandSimRequestWrapper.portalIfc;
   portals[1] = nandSimIndicationProxy.portalIfc; 

   portals[2] = strstrRequestWrapper.portalIfc;
   portals[3] = strstrIndicationProxy.portalIfc; 
   
   portals[4] = backingStoreSGListConfigRequestWrapper.portalIfc;
   portals[5] = backingStoreSGListConfigIndicationProxy.portalIfc;

   portals[6] = nandsimSGListConfigRequestWrapper.portalIfc;
   portals[7] = nandsimSGListConfigIndicationProxy.portalIfc;
   
   portals[8] = hostDmaDebugRequestWrapper.portalIfc;
   portals[9] = hostDmaDebugIndicationProxy.portalIfc; 

   portals[10] = nandsimDmaRequestWrapper.portalIfc;
   portals[11] = nandsimDmaDebugIndicationProxy.portalIfc; 
   
   portals[12] = algoSGListConfigRequestWrapper.portalIfc;
   portals[13] = algoSGListConfigIndicationProxy.portalIfc;

   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = hostDma.masters;
   interface leds = default_leds;
      
endmodule : mkPortalTop
