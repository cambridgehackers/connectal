
// Copyright (c) 2013 Quanta Research Cambridge, Inc.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

import Clocks       :: *;
import DefaultValue :: *;
import XilinxCells  :: *;
import Vector       :: *;

(* always_ready, always_enabled *)
interface Ps7#(numeric type C_EMIO_GPIO_WIDTH);
    method Action CAN0_PHY_RX(Bit#(1) v);
    method Bit#(1) CAN0_PHY_TX();
    method Action CAN1_PHY_RX(Bit#(1) v);
    method Bit#(1) CAN1_PHY_TX();
    method Action Core0_nFIQ(Bit#(1) v);
    method Action Core0_nIRQ(Bit#(1) v);
    method Action Core1_nFIQ(Bit#(1) v);
    method Action Core1_nIRQ(Bit#(1) v);
    method Action DDR_ARB(Bit#(4) v);
    method Bit#(15) DDR_Addr();
    method Bit#(3) DDR_BankAddr();
    method Bit#(1) DDR_CAS_n();
    method Bit#(1) DDR_CKE();
    method Bit#(1) DDR_CS_n();
    method Bit#(1) DDR_Clk();
    method Bit#(1) DDR_Clk_n();
    method Bit#(C_DM_WIDTH) DDR_DM();
    method Bit#(C_DQ_WIDTH) DDR_DQ();
    method Bit#(C_DQS_WIDTH) DDR_DQS();
    method Bit#(C_DQS_WIDTH) DDR_DQS_n();
    method Bit#(1) DDR_DRSTB();
    method Bit#(1) DDR_ODT();
    method Bit#(1) DDR_RAS_n();
    method Bit#(1) DDR_VRN();
    method Bit#(1) DDR_VRP();
    method Bit#(1) DDR_WEB();
    method Action DMA0_ACLK(Bit#(1) v);
    method Action DMA0_DAREADY(Bit#(1) v);
    method Bit#(2) DMA0_DATYPE();
    method Bit#(1) DMA0_DAVALID();
    method Action DMA0_DRLAST(Bit#(1) v);
    method Bit#(1) DMA0_DRREADY();
    method Action DMA0_DRTYPE(Bit#(2) v);
    method Action DMA0_DRVALID(Bit#(1) v);
    method Bit#(1) DMA0_RSTN();
    method Action DMA1_ACLK(Bit#(1) v);
    method Action DMA1_DAREADY(Bit#(1) v);
    method Bit#(2) DMA1_DATYPE();
    method Bit#(1) DMA1_DAVALID();
    method Action DMA1_DRLAST(Bit#(1) v);
    method Bit#(1) DMA1_DRREADY();
    method Action DMA1_DRTYPE(Bit#(2) v);
    method Action DMA1_DRVALID(Bit#(1) v);
    method Bit#(1) DMA1_RSTN();
    method Action DMA2_ACLK(Bit#(1) v);
    method Action DMA2_DAREADY(Bit#(1) v);
    method Bit#(2) DMA2_DATYPE();
    method Bit#(1) DMA2_DAVALID();
    method Action DMA2_DRLAST(Bit#(1) v);
    method Bit#(1) DMA2_DRREADY();
    method Action DMA2_DRTYPE(Bit#(2) v);
    method Action DMA2_DRVALID(Bit#(1) v);
    method Bit#(1) DMA2_RSTN();
    method Action DMA3_ACLK(Bit#(1) v);
    method Action DMA3_DAREADY(Bit#(1) v);
    method Bit#(2) DMA3_DATYPE();
    method Bit#(1) DMA3_DAVALID();
    method Action DMA3_DRLAST(Bit#(1) v);
    method Bit#(1) DMA3_DRREADY();
    method Action DMA3_DRTYPE(Bit#(2) v);
    method Action DMA3_DRVALID(Bit#(1) v);
    method Bit#(1) DMA3_RSTN();
    method Action ENET0_EXT_INTIN(Bit#(1) v);
    method Action ENET0_GMII_COL(Bit#(1) v);
    method Action ENET0_GMII_CRS(Bit#(1) v);
    method Action ENET0_GMII_RXD(Bit#(8) v);
    method Action ENET0_GMII_RX_CLK(Bit#(1) v);
    method Action ENET0_GMII_RX_DV(Bit#(1) v);
    method Action ENET0_GMII_RX_ER(Bit#(1) v);
    method Bit#(8) ENET0_GMII_TXD();
    method Action ENET0_GMII_TX_CLK(Bit#(1) v);
    method Bit#(1) ENET0_GMII_TX_EN();
    method Bit#(1) ENET0_GMII_TX_ER();
    method Action ENET0_MDIO_I(Bit#(1) v);
    method Bit#(1) ENET0_MDIO_MDC();
    method Bit#(1) ENET0_MDIO_O();
    method Bit#(1) ENET0_MDIO_T();
    method Bit#(1) ENET0_PTP_DELAY_REQ_RX();
    method Bit#(1) ENET0_PTP_DELAY_REQ_TX();
    method Bit#(1) ENET0_PTP_PDELAY_REQ_RX();
    method Bit#(1) ENET0_PTP_PDELAY_REQ_TX();
    method Bit#(1) ENET0_PTP_PDELAY_RESP_RX();
    method Bit#(1) ENET0_PTP_PDELAY_RESP_TX();
    method Bit#(1) ENET0_PTP_SYNC_FRAME_RX();
    method Bit#(1) ENET0_PTP_SYNC_FRAME_TX();
    method Bit#(1) ENET0_SOF_RX();
    method Bit#(1) ENET0_SOF_TX();
    method Action ENET1_EXT_INTIN(Bit#(1) v);
    method Action ENET1_GMII_COL(Bit#(1) v);
    method Action ENET1_GMII_CRS(Bit#(1) v);
    method Action ENET1_GMII_RXD(Bit#(8) v);
    method Action ENET1_GMII_RX_CLK(Bit#(1) v);
    method Action ENET1_GMII_RX_DV(Bit#(1) v);
    method Action ENET1_GMII_RX_ER(Bit#(1) v);
    method Bit#(8) ENET1_GMII_TXD();
    method Action ENET1_GMII_TX_CLK(Bit#(1) v);
    method Bit#(1) ENET1_GMII_TX_EN();
    method Bit#(1) ENET1_GMII_TX_ER();
    method Action ENET1_MDIO_I(Bit#(1) v);
    method Bit#(1) ENET1_MDIO_MDC();
    method Bit#(1) ENET1_MDIO_O();
    method Bit#(1) ENET1_MDIO_T();
    method Bit#(1) ENET1_PTP_DELAY_REQ_RX();
    method Bit#(1) ENET1_PTP_DELAY_REQ_TX();
    method Bit#(1) ENET1_PTP_PDELAY_REQ_RX();
    method Bit#(1) ENET1_PTP_PDELAY_REQ_TX();
    method Bit#(1) ENET1_PTP_PDELAY_RESP_RX();
    method Bit#(1) ENET1_PTP_PDELAY_RESP_TX();
    method Bit#(1) ENET1_PTP_SYNC_FRAME_RX();
    method Bit#(1) ENET1_PTP_SYNC_FRAME_TX();
    method Bit#(1) ENET1_SOF_RX();
    method Bit#(1) ENET1_SOF_TX();
    method Action EVENT_EVENTI(Bit#(1) v);
    method Bit#(1) EVENT_EVENTO();
    method Bit#(2) EVENT_STANDBYWFE();
    method Bit#(2) EVENT_STANDBYWFI();
    method Bit#(1) FCLK_CLK0();
    method Bit#(1) FCLK_CLK1();
    method Bit#(1) FCLK_CLK2();
    method Bit#(1) FCLK_CLK3();
    method Action FCLK_CLKTRIG0_N(Bit#(1) v);
    method Action FCLK_CLKTRIG1_N(Bit#(1) v);
    method Action FCLK_CLKTRIG2_N(Bit#(1) v);
    method Action FCLK_CLKTRIG3_N(Bit#(1) v);
    method Bit#(1) FCLK_RESET0_N();
    method Bit#(1) FCLK_RESET1_N();
    method Bit#(1) FCLK_RESET2_N();
    method Bit#(1) FCLK_RESET3_N();
    method Action FPGA_IDLE_N(Bit#(1) v);
    method Action FTMD_TRACEIN_ATID(Bit#(4) v);
    method Action FTMD_TRACEIN_CLK(Bit#(1) v);
    method Action FTMD_TRACEIN_DATA(Bit#(32) v);
    method Action FTMD_TRACEIN_VALID(Bit#(1) v);
    method Action FTMT_F2P_DEBUG(Bit#(32) v);
    method Action FTMT_F2P_TRIG(Bit#(4) v);
    method Bit#(4) FTMT_F2P_TRIGACK();
    method Bit#(32) FTMT_P2F_DEBUG();
    method Bit#(4) FTMT_P2F_TRIG();
    method Action FTMT_P2F_TRIGACK(Bit#(4) v);
    method Action GPIO_I(Bit#(C_EMIO_GPIO_WIDTH) v);
    method Bit#(C_EMIO_GPIO_WIDTH) GPIO_O();
    method Bit#(C_EMIO_GPIO_WIDTH) GPIO_T();
    method Action I2C0_SCL_I(Bit#(1) v);
    method Bit#(1) I2C0_SCL_O();
    method Bit#(1) I2C0_SCL_T();
    method Action I2C0_SDA_I(Bit#(1) v);
    method Bit#(1) I2C0_SDA_O();
    method Bit#(1) I2C0_SDA_T();
    method Action I2C1_SCL_I(Bit#(1) v);
    method Bit#(1) I2C1_SCL_O();
    method Bit#(1) I2C1_SCL_T();
    method Action I2C1_SDA_I(Bit#(1) v);
    method Bit#(1) I2C1_SDA_O();
    method Bit#(1) I2C1_SDA_T();
    method Action IRQ_F2P(Bit#(16) v);
    method Bit#(1) IRQ_P2F_CAN0();
    method Bit#(1) IRQ_P2F_CAN1();
    method Bit#(1) IRQ_P2F_CTI();
    method Bit#(1) IRQ_P2F_DMAC0();
    method Bit#(1) IRQ_P2F_DMAC1();
    method Bit#(1) IRQ_P2F_DMAC2();
    method Bit#(1) IRQ_P2F_DMAC3();
    method Bit#(1) IRQ_P2F_DMAC4();
    method Bit#(1) IRQ_P2F_DMAC5();
    method Bit#(1) IRQ_P2F_DMAC6();
    method Bit#(1) IRQ_P2F_DMAC7();
    method Bit#(1) IRQ_P2F_DMAC_ABORT();
    method Bit#(1) IRQ_P2F_ENET0();
    method Bit#(1) IRQ_P2F_ENET1();
    method Bit#(1) IRQ_P2F_ENET_WAKE0();
    method Bit#(1) IRQ_P2F_ENET_WAKE1();
    method Bit#(1) IRQ_P2F_GPIO();
    method Bit#(1) IRQ_P2F_I2C0();
    method Bit#(1) IRQ_P2F_I2C1();
    method Bit#(1) IRQ_P2F_QSPI();
    method Bit#(1) IRQ_P2F_SDIO0();
    method Bit#(1) IRQ_P2F_SDIO1();
    method Bit#(1) IRQ_P2F_SMC();
    method Bit#(1) IRQ_P2F_SPI0();
    method Bit#(1) IRQ_P2F_SPI1();
    method Bit#(1) IRQ_P2F_UART0();
    method Bit#(1) IRQ_P2F_UART1();
    method Bit#(1) IRQ_P2F_USB0();
    method Bit#(1) IRQ_P2F_USB1();
    method Bit#(C_MIO_PRIMITIVE) MIO();
    method Action M_AXI_GP0_ACLK(Bit#(1) v);
    method Bit#(32) M_AXI_GP0_ARADDR();
    method Bit#(2) M_AXI_GP0_ARBURST();
    method Bit#(4) M_AXI_GP0_ARCACHE();
    method Bit#(1) M_AXI_GP0_ARESETN();
    method Bit#(C_M_AXI_GP0_THREAD_ID_WIDTH) M_AXI_GP0_ARID();
    method Bit#(4) M_AXI_GP0_ARLEN();
    method Bit#(2) M_AXI_GP0_ARLOCK();
    method Bit#(3) M_AXI_GP0_ARPROT();
    method Bit#(4) M_AXI_GP0_ARQOS();
    method Action M_AXI_GP0_ARREADY(Bit#(1) v);
    method Bit#(3) M_AXI_GP0_ARSIZE();
    method Bit#(1) M_AXI_GP0_ARVALID();
    method Bit#(32) M_AXI_GP0_AWADDR();
    method Bit#(2) M_AXI_GP0_AWBURST();
    method Bit#(4) M_AXI_GP0_AWCACHE();
    method Bit#(C_M_AXI_GP0_THREAD_ID_WIDTH) M_AXI_GP0_AWID();
    method Bit#(4) M_AXI_GP0_AWLEN();
    method Bit#(2) M_AXI_GP0_AWLOCK();
    method Bit#(3) M_AXI_GP0_AWPROT();
    method Bit#(4) M_AXI_GP0_AWQOS();
    method Action M_AXI_GP0_AWREADY(Bit#(1) v);
    method Bit#(3) M_AXI_GP0_AWSIZE();
    method Bit#(1) M_AXI_GP0_AWVALID();
    method Action M_AXI_GP0_BID(Bit#(C_M_AXI_GP0_THREAD_ID_WIDTH) v);
    method Bit#(1) M_AXI_GP0_BREADY();
    method Action M_AXI_GP0_BRESP(Bit#(2) v);
    method Action M_AXI_GP0_BVALID(Bit#(1) v);
    method Action M_AXI_GP0_RDATA(Bit#(32) v);
    method Action M_AXI_GP0_RID(Bit#(C_M_AXI_GP0_THREAD_ID_WIDTH) v);
    method Action M_AXI_GP0_RLAST(Bit#(1) v);
    method Bit#(1) M_AXI_GP0_RREADY();
    method Action M_AXI_GP0_RRESP(Bit#(2) v);
    method Action M_AXI_GP0_RVALID(Bit#(1) v);
    method Bit#(32) M_AXI_GP0_WDATA();
    method Bit#(C_M_AXI_GP0_THREAD_ID_WIDTH) M_AXI_GP0_WID();
    method Bit#(1) M_AXI_GP0_WLAST();
    method Action M_AXI_GP0_WREADY(Bit#(1) v);
    method Bit#(4) M_AXI_GP0_WSTRB();
    method Bit#(1) M_AXI_GP0_WVALID();
    method Action M_AXI_GP1_ACLK(Bit#(1) v);
    method Bit#(32) M_AXI_GP1_ARADDR();
    method Bit#(2) M_AXI_GP1_ARBURST();
    method Bit#(4) M_AXI_GP1_ARCACHE();
    method Bit#(1) M_AXI_GP1_ARESETN();
    method Bit#(C_M_AXI_GP1_THREAD_ID_WIDTH) M_AXI_GP1_ARID();
    method Bit#(4) M_AXI_GP1_ARLEN();
    method Bit#(2) M_AXI_GP1_ARLOCK();
    method Bit#(3) M_AXI_GP1_ARPROT();
    method Bit#(4) M_AXI_GP1_ARQOS();
    method Action M_AXI_GP1_ARREADY(Bit#(1) v);
    method Bit#(3) M_AXI_GP1_ARSIZE();
    method Bit#(1) M_AXI_GP1_ARVALID();
    method Bit#(32) M_AXI_GP1_AWADDR();
    method Bit#(2) M_AXI_GP1_AWBURST();
    method Bit#(4) M_AXI_GP1_AWCACHE();
    method Bit#(C_M_AXI_GP1_THREAD_ID_WIDTH) M_AXI_GP1_AWID();
    method Bit#(4) M_AXI_GP1_AWLEN();
    method Bit#(2) M_AXI_GP1_AWLOCK();
    method Bit#(3) M_AXI_GP1_AWPROT();
    method Bit#(4) M_AXI_GP1_AWQOS();
    method Action M_AXI_GP1_AWREADY(Bit#(1) v);
    method Bit#(3) M_AXI_GP1_AWSIZE();
    method Bit#(1) M_AXI_GP1_AWVALID();
    method Action M_AXI_GP1_BID(Bit#(C_M_AXI_GP1_THREAD_ID_WIDTH) v);
    method Bit#(1) M_AXI_GP1_BREADY();
    method Action M_AXI_GP2_BRESP(Bit#(1) v);
    method Action M_AXI_GP1_BVALID(Bit#(1) v);
    method Action M_AXI_GP1_RDATA(Bit#(32) v);
    method Action M_AXI_GP1_RID(Bit#(C_M_AXI_GP1_THREAD_ID_WIDTH) v);
    method Action M_AXI_GP1_RLAST(Bit#(1) v);
    method Bit#(1) M_AXI_GP1_RREADY();
    method Action M_AXI_GP2_RRESP(Bit#(1) v);
    method Action M_AXI_GP1_RVALID(Bit#(1) v);
    method Bit#(32) M_AXI_GP1_WDATA();
    method Bit#(C_M_AXI_GP1_THREAD_ID_WIDTH) M_AXI_GP1_WID();
    method Bit#(1) M_AXI_GP1_WLAST();
    method Action M_AXI_GP1_WREADY(Bit#(1) v);
    method Bit#(4) M_AXI_GP1_WSTRB();
    method Bit#(1) M_AXI_GP1_WVALID();
    method Action PJTAG_TCK(Bit#(1) v);
    method Action PJTAG_TD_I(Bit#(1) v);
    method Bit#(1) PJTAG_TD_O();
    method Bit#(1) PJTAG_TD_T();
    method Action PJTAG_TMS(Bit#(1) v);
    method Action PS_CLK(Bit#(1) v);
    method Action PS_PORB(Bit#(1) v);
    method Action PS_SRSTB(Bit#(1) v);
    method Bit#(1) SDIO0_BUSPOW();
    method Bit#(3) SDIO0_BUSVOLT();
    method Action SDIO0_CDN(Bit#(1) v);
    method Bit#(1) SDIO0_CLK();
    method Action SDIO0_CLK_FB(Bit#(1) v);
    method Action SDIO0_CMD_I(Bit#(1) v);
    method Bit#(1) SDIO0_CMD_O();
    method Bit#(1) SDIO0_CMD_T();
    method Action SDIO0_DATA_I(Bit#(4) v);
    method Bit#(4) SDIO0_DATA_O();
    method Bit#(4) SDIO0_DATA_T();
    method Bit#(1) SDIO0_LED();
    method Action SDIO0_WP(Bit#(1) v);
    method Bit#(1) SDIO1_BUSPOW();
    method Bit#(3) SDIO1_BUSVOLT();
    method Action SDIO1_CDN(Bit#(1) v);
    method Bit#(1) SDIO1_CLK();
    method Action SDIO1_CLK_FB(Bit#(1) v);
    method Action SDIO1_CMD_I(Bit#(1) v);
    method Bit#(1) SDIO1_CMD_O();
    method Bit#(1) SDIO1_CMD_T();
    method Action SDIO1_DATA_I(Bit#(4) v);
    method Bit#(4) SDIO1_DATA_O();
    method Bit#(4) SDIO1_DATA_T();
    method Bit#(1) SDIO1_LED();
    method Action SDIO1_WP(Bit#(1) v);
    method Action SPI0_MISO_I(Bit#(1) v);
    method Bit#(1) SPI0_MISO_O();
    method Bit#(1) SPI0_MISO_T();
    method Action SPI0_MOSI_I(Bit#(1) v);
    method Bit#(1) SPI0_MOSI_O();
    method Bit#(1) SPI0_MOSI_T();
    method Action SPI0_SCLK_I(Bit#(1) v);
    method Bit#(1) SPI0_SCLK_O();
    method Bit#(1) SPI0_SCLK_T();
    method Bit#(1) SPI0_SS1_O();
    method Bit#(1) SPI0_SS2_O();
    method Action SPI0_SS_I(Bit#(1) v);
    method Bit#(1) SPI0_SS_O();
    method Bit#(1) SPI0_SS_T();
    method Action SPI1_MISO_I(Bit#(1) v);
    method Bit#(1) SPI1_MISO_O();
    method Bit#(1) SPI1_MISO_T();
    method Action SPI1_MOSI_I(Bit#(1) v);
    method Bit#(1) SPI1_MOSI_O();
    method Bit#(1) SPI1_MOSI_T();
    method Action SPI1_SCLK_I(Bit#(1) v);
    method Bit#(1) SPI1_SCLK_O();
    method Bit#(1) SPI1_SCLK_T();
    method Bit#(1) SPI1_SS1_O();
    method Bit#(1) SPI1_SS2_O();
    method Action SPI1_SS_I(Bit#(1) v);
    method Bit#(1) SPI1_SS_O();
    method Bit#(1) SPI1_SS_T();
    method Action SRAM_INTIN(Bit#(1) v);
    method Action S_AXI_ACP_ACLK(Bit#(1) v);
    method Action S_AXI_ACP_ARADDR(Bit#(32) v);
    method Action S_AXI_ACP_ARBURST(Bit#(2) v);
    method Action S_AXI_ACP_ARCACHE(Bit#(4) v);
    method Bit#(1) S_AXI_ACP_ARESETN();
    method Action S_AXI_ACP_ARID(Bit#(C_S_AXI_ACP_ID_WIDTH) v);
    method Action S_AXI_ACP_ARLEN(Bit#(4) v);
    method Action S_AXI_ACP_ARLOCK(Bit#(2) v);
    method Action S_AXI_ACP_ARPROT(Bit#(3) v);
    method Action S_AXI_ACP_ARQOS(Bit#(4) v);
    method Bit#(1) S_AXI_ACP_ARREADY();
    method Action S_AXI_ACP_ARSIZE(Bit#(3) v);
    method Action S_AXI_ACP_ARUSER(Bit#(5) v);
    method Action S_AXI_ACP_ARVALID(Bit#(1) v);
    method Action S_AXI_ACP_AWADDR(Bit#(32) v);
    method Action S_AXI_ACP_AWBURST(Bit#(2) v);
    method Action S_AXI_ACP_AWCACHE(Bit#(4) v);
    method Action S_AXI_ACP_AWID(Bit#(C_S_AXI_ACP_ID_WIDTH) v);
    method Action S_AXI_ACP_AWLEN(Bit#(4) v);
    method Action S_AXI_ACP_AWLOCK(Bit#(2) v);
    method Action S_AXI_ACP_AWPROT(Bit#(3) v);
    method Action S_AXI_ACP_AWQOS(Bit#(4) v);
    method Bit#(1) S_AXI_ACP_AWREADY();
    method Action S_AXI_ACP_AWSIZE(Bit#(3) v);
    method Action S_AXI_ACP_AWUSER(Bit#(5) v);
    method Action S_AXI_ACP_AWVALID(Bit#(1) v);
    method Bit#(C_S_AXI_ACP_ID_WIDTH) S_AXI_ACP_BID();
    method Action S_AXI_ACP_BREADY(Bit#(1) v);
    method Bit#(2) S_AXI_ACP_BRESP();
    method Bit#(1) S_AXI_ACP_BVALID();
    method Bit#(64) S_AXI_ACP_RDATA();
    method Bit#(C_S_AXI_ACP_ID_WIDTH) S_AXI_ACP_RID();
    method Bit#(1) S_AXI_ACP_RLAST();
    method Action S_AXI_ACP_RREADY(Bit#(1) v);
    method Bit#(2) S_AXI_ACP_RRESP();
    method Bit#(1) S_AXI_ACP_RVALID();
    method Action S_AXI_ACP_WDATA(Bit#(64) v);
    method Action S_AXI_ACP_WID(Bit#(C_S_AXI_ACP_ID_WIDTH) v);
    method Action S_AXI_ACP_WLAST(Bit#(1) v);
    method Bit#(1) S_AXI_ACP_WREADY();
    method Action S_AXI_ACP_WSTRB(Bit#(8) v);
    method Action S_AXI_ACP_WVALID(Bit#(1) v);
    method Action S_AXI_GP0_ACLK(Bit#(1) v);
    method Action S_AXI_GP0_ARADDR(Bit#(32) v);
    method Action S_AXI_GP0_ARBURST(Bit#(2) v);
    method Action S_AXI_GP0_ARCACHE(Bit#(4) v);
    method Bit#(1) S_AXI_GP0_ARESETN();
    method Action S_AXI_GP0_ARID(Bit#(C_S_AXI_GP0_ID_WIDTH) v);
    method Action S_AXI_GP0_ARLEN(Bit#(4) v);
    method Action S_AXI_GP0_ARLOCK(Bit#(2) v);
    method Action S_AXI_GP0_ARPROT(Bit#(3) v);
    method Action S_AXI_GP0_ARQOS(Bit#(4) v);
    method Bit#(1) S_AXI_GP0_ARREADY();
    method Action S_AXI_GP0_ARSIZE(Bit#(3) v);
    method Action S_AXI_GP0_ARVALID(Bit#(1) v);
    method Action S_AXI_GP0_AWADDR(Bit#(32) v);
    method Action S_AXI_GP0_AWBURST(Bit#(2) v);
    method Action S_AXI_GP0_AWCACHE(Bit#(4) v);
    method Action S_AXI_GP0_AWID(Bit#(C_S_AXI_GP0_ID_WIDTH) v);
    method Action S_AXI_GP0_AWLEN(Bit#(4) v);
    method Action S_AXI_GP0_AWLOCK(Bit#(2) v);
    method Action S_AXI_GP0_AWPROT(Bit#(3) v);
    method Action S_AXI_GP0_AWQOS(Bit#(4) v);
    method Bit#(1) S_AXI_GP0_AWREADY();
    method Action S_AXI_GP0_AWSIZE(Bit#(3) v);
    method Action S_AXI_GP0_AWVALID(Bit#(1) v);
    method Bit#(C_S_AXI_GP0_ID_WIDTH) S_AXI_GP0_BID();
    method Action S_AXI_GP0_BREADY(Bit#(1) v);
    method Bit#(2) S_AXI_GP0_BRESP();
    method Bit#(1) S_AXI_GP0_BVALID();
    method Bit#(32) S_AXI_GP0_RDATA();
    method Bit#(C_S_AXI_GP0_ID_WIDTH) S_AXI_GP0_RID();
    method Bit#(1) S_AXI_GP0_RLAST();
    method Action S_AXI_GP0_RREADY(Bit#(1) v);
    method Bit#(2) S_AXI_GP0_RRESP();
    method Bit#(1) S_AXI_GP0_RVALID();
    method Action S_AXI_GP0_WDATA(Bit#(32) v);
    method Action S_AXI_GP0_WID(Bit#(C_S_AXI_GP0_ID_WIDTH) v);
    method Action S_AXI_GP0_WLAST(Bit#(1) v);
    method Bit#(1) S_AXI_GP0_WREADY();
    method Action S_AXI_GP0_WSTRB(Bit#(4) v);
    method Action S_AXI_GP0_WVALID(Bit#(1) v);
    method Action S_AXI_GP1_ACLK(Bit#(1) v);
    method Action S_AXI_GP1_ARADDR(Bit#(32) v);
    method Action S_AXI_GP2_ARBURST(Bit#(1) v);
    method Action S_AXI_GP1_ARCACHE(Bit#(4) v);
    method Bit#(1) S_AXI_GP1_ARESETN();
    method Action S_AXI_GP1_ARID(Bit#(C_S_AXI_GP1_ID_WIDTH) v);
    method Action S_AXI_GP1_ARLEN(Bit#(4) v);
    method Action S_AXI_GP2_ARLOCK(Bit#(1) v);
    method Action S_AXI_GP1_ARPROT(Bit#(3) v);
    method Action S_AXI_GP1_ARQOS(Bit#(4) v);
    method Bit#(1) S_AXI_GP1_ARREADY();
    method Action S_AXI_GP1_ARSIZE(Bit#(3) v);
    method Action S_AXI_GP1_ARVALID(Bit#(1) v);
    method Action S_AXI_GP1_AWADDR(Bit#(32) v);
    method Action S_AXI_GP2_AWBURST(Bit#(1) v);
    method Action S_AXI_GP1_AWCACHE(Bit#(4) v);
    method Action S_AXI_GP1_AWID(Bit#(C_S_AXI_GP1_ID_WIDTH) v);
    method Action S_AXI_GP1_AWLEN(Bit#(4) v);
    method Action S_AXI_GP2_AWLOCK(Bit#(1) v);
    method Action S_AXI_GP1_AWPROT(Bit#(3) v);
    method Action S_AXI_GP1_AWQOS(Bit#(4) v);
    method Bit#(1) S_AXI_GP1_AWREADY();
    method Action S_AXI_GP1_AWSIZE(Bit#(3) v);
    method Action S_AXI_GP1_AWVALID(Bit#(1) v);
    method Bit#(C_S_AXI_GP1_ID_WIDTH) S_AXI_GP1_BID();
    method Action S_AXI_GP1_BREADY(Bit#(1) v);
    method Bit#(2) S_AXI_GP1_BRESP();
    method Bit#(1) S_AXI_GP1_BVALID();
    method Bit#(32) S_AXI_GP1_RDATA();
    method Bit#(C_S_AXI_GP1_ID_WIDTH) S_AXI_GP1_RID();
    method Bit#(1) S_AXI_GP1_RLAST();
    method Action S_AXI_GP1_RREADY(Bit#(1) v);
    method Bit#(2) S_AXI_GP1_RRESP();
    method Bit#(1) S_AXI_GP1_RVALID();
    method Action S_AXI_GP1_WDATA(Bit#(32) v);
    method Action S_AXI_GP1_WID(Bit#(C_S_AXI_GP1_ID_WIDTH) v);
    method Action S_AXI_GP1_WLAST(Bit#(1) v);
    method Bit#(1) S_AXI_GP1_WREADY();
    method Action S_AXI_GP1_WSTRB(Bit#(4) v);
    method Action S_AXI_GP1_WVALID(Bit#(1) v);
    method Action S_AXI_HP0_ACLK(Bit#(1) v);
    method Action S_AXI_HP0_ARADDR(Bit#(32) v);
    method Action S_AXI_HP0_ARBURST(Bit#(2) v);
    method Action S_AXI_HP0_ARCACHE(Bit#(4) v);
    method Bit#(1) S_AXI_HP0_ARESETN();
    method Action S_AXI_HP0_ARID(Bit#(C_S_AXI_HP0_ID_WIDTH) v);
    method Action S_AXI_HP0_ARLEN(Bit#(4) v);
    method Action S_AXI_HP0_ARLOCK(Bit#(2) v);
    method Action S_AXI_HP0_ARPROT(Bit#(3) v);
    method Action S_AXI_HP0_ARQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP0_ARREADY();
    method Action S_AXI_HP0_ARSIZE(Bit#(3) v);
    method Action S_AXI_HP0_ARVALID(Bit#(1) v);
    method Action S_AXI_HP0_AWADDR(Bit#(32) v);
    method Action S_AXI_HP0_AWBURST(Bit#(2) v);
    method Action S_AXI_HP0_AWCACHE(Bit#(4) v);
    method Action S_AXI_HP0_AWID(Bit#(C_S_AXI_HP0_ID_WIDTH) v);
    method Action S_AXI_HP0_AWLEN(Bit#(4) v);
    method Action S_AXI_HP0_AWLOCK(Bit#(2) v);
    method Action S_AXI_HP0_AWPROT(Bit#(3) v);
    method Action S_AXI_HP0_AWQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP0_AWREADY();
    method Action S_AXI_HP0_AWSIZE(Bit#(3) v);
    method Action S_AXI_HP0_AWVALID(Bit#(1) v);
    method Bit#(C_S_AXI_HP0_ID_WIDTH) S_AXI_HP0_BID();
    method Action S_AXI_HP0_BREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP0_BRESP();
    method Bit#(1) S_AXI_HP0_BVALID();
    method Bit#(3) S_AXI_HP0_RACOUNT();
    method Bit#(8) S_AXI_HP0_RCOUNT();
    method Bit#(C_S_AXI_HP0_DATA_WIDTH) S_AXI_HP0_RDATA();
    method Action S_AXI_HP0_RDISSUECAP1_EN(Bit#(1) v);
    method Bit#(C_S_AXI_HP0_ID_WIDTH) S_AXI_HP0_RID();
    method Bit#(1) S_AXI_HP0_RLAST();
    method Action S_AXI_HP0_RREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP0_RRESP();
    method Bit#(1) S_AXI_HP0_RVALID();
    method Bit#(6) S_AXI_HP0_WACOUNT();
    method Bit#(8) S_AXI_HP0_WCOUNT();
    method Action S_AXI_HP0_WDATA(Bit#(C_S_AXI_HP0_DATA_WIDTH) v);
    method Action S_AXI_HP0_WID(Bit#(C_S_AXI_HP0_ID_WIDTH) v);
    method Action S_AXI_HP0_WLAST(Bit#(1) v);
    method Bit#(1) S_AXI_HP0_WREADY();
    method Action S_AXI_HP0_WRISSUECAP1_EN(Bit#(1) v);
    method Action S_AXI_HP0_WSTRB(Bit#(C_S_AXI_HP0_DATA_WIDTH/8) v);
    method Action S_AXI_HP0_WVALID(Bit#(1) v);
    method Action S_AXI_HP1_ACLK(Bit#(1) v);
    method Action S_AXI_HP1_ARADDR(Bit#(32) v);
    method Action S_AXI_HP2_ARBURST(Bit#(1) v);
    method Action S_AXI_HP1_ARCACHE(Bit#(4) v);
    method Bit#(1) S_AXI_HP1_ARESETN();
    method Action S_AXI_HP1_ARID(Bit#(C_S_AXI_HP1_ID_WIDTH) v);
    method Action S_AXI_HP1_ARLEN(Bit#(4) v);
    method Action S_AXI_HP2_ARLOCK(Bit#(1) v);
    method Action S_AXI_HP1_ARPROT(Bit#(3) v);
    method Action S_AXI_HP1_ARQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP1_ARREADY();
    method Action S_AXI_HP1_ARSIZE(Bit#(3) v);
    method Action S_AXI_HP1_ARVALID(Bit#(1) v);
    method Action S_AXI_HP1_AWADDR(Bit#(32) v);
    method Action S_AXI_HP2_AWBURST(Bit#(1) v);
    method Action S_AXI_HP1_AWCACHE(Bit#(4) v);
    method Action S_AXI_HP1_AWID(Bit#(C_S_AXI_HP1_ID_WIDTH) v);
    method Action S_AXI_HP1_AWLEN(Bit#(4) v);
    method Action S_AXI_HP2_AWLOCK(Bit#(1) v);
    method Action S_AXI_HP1_AWPROT(Bit#(3) v);
    method Action S_AXI_HP1_AWQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP1_AWREADY();
    method Action S_AXI_HP1_AWSIZE(Bit#(3) v);
    method Action S_AXI_HP1_AWVALID(Bit#(1) v);
    method Bit#(C_S_AXI_HP1_ID_WIDTH) S_AXI_HP1_BID();
    method Action S_AXI_HP1_BREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP1_BRESP();
    method Bit#(1) S_AXI_HP1_BVALID();
    method Bit#(3) S_AXI_HP1_RACOUNT();
    method Bit#(8) S_AXI_HP1_RCOUNT();
    method Bit#(C_S_AXI_HP1_DATA_WIDTH) S_AXI_HP1_RDATA();
    method Action S_AXI_HP1_RDISSUECAP1_EN(Bit#(1) v);
    method Bit#(C_S_AXI_HP1_ID_WIDTH) S_AXI_HP1_RID();
    method Bit#(1) S_AXI_HP1_RLAST();
    method Action S_AXI_HP1_RREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP1_RRESP();
    method Bit#(1) S_AXI_HP1_RVALID();
    method Bit#(6) S_AXI_HP1_WACOUNT();
    method Bit#(8) S_AXI_HP1_WCOUNT();
    method Action S_AXI_HP1_WDATA(Bit#(C_S_AXI_HP1_DATA_WIDTH) v);
    method Action S_AXI_HP1_WID(Bit#(C_S_AXI_HP1_ID_WIDTH) v);
    method Action S_AXI_HP1_WLAST(Bit#(1) v);
    method Bit#(1) S_AXI_HP1_WREADY();
    method Action S_AXI_HP1_WRISSUECAP1_EN(Bit#(1) v);
    method Action S_AXI_HP1_WSTRB(Bit#(C_S_AXI_HP1_DATA_WIDTH) v);
    method Action S_AXI_HP1_WVALID(Bit#(1) v);
    method Action S_AXI_HP2_ACLK(Bit#(1) v);
    method Action S_AXI_HP2_ARADDR(Bit#(32) v);
    method Action S_AXI_HP2_ARBURST(Bit#(2) v);
    method Action S_AXI_HP2_ARCACHE(Bit#(4) v);
    method Bit#(1) S_AXI_HP2_ARESETN();
    method Action S_AXI_HP2_ARID(Bit#(C_S_AXI_HP2_ID_WIDTH) v);
    method Action S_AXI_HP2_ARLEN(Bit#(4) v);
    method Action S_AXI_HP2_ARLOCK(Bit#(2) v);
    method Action S_AXI_HP2_ARPROT(Bit#(3) v);
    method Action S_AXI_HP2_ARQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP2_ARREADY();
    method Action S_AXI_HP2_ARSIZE(Bit#(3) v);
    method Action S_AXI_HP2_ARVALID(Bit#(1) v);
    method Action S_AXI_HP2_AWADDR(Bit#(32) v);
    method Action S_AXI_HP2_AWBURST(Bit#(2) v);
    method Action S_AXI_HP2_AWCACHE(Bit#(4) v);
    method Action S_AXI_HP2_AWID(Bit#(C_S_AXI_HP2_ID_WIDTH) v);
    method Action S_AXI_HP2_AWLEN(Bit#(4) v);
    method Action S_AXI_HP2_AWLOCK(Bit#(2) v);
    method Action S_AXI_HP2_AWPROT(Bit#(3) v);
    method Action S_AXI_HP2_AWQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP2_AWREADY();
    method Action S_AXI_HP2_AWSIZE(Bit#(3) v);
    method Action S_AXI_HP2_AWVALID(Bit#(1) v);
    method Bit#(C_S_AXI_HP2_ID_WIDTH) S_AXI_HP2_BID();
    method Action S_AXI_HP2_BREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP2_BRESP();
    method Bit#(1) S_AXI_HP2_BVALID();
    method Bit#(3) S_AXI_HP2_RACOUNT();
    method Bit#(8) S_AXI_HP2_RCOUNT();
    method Bit#(C_S_AXI_HP2_DATA_WIDTH) S_AXI_HP2_RDATA();
    method Action S_AXI_HP2_RDISSUECAP1_EN(Bit#(1) v);
    method Bit#(C_S_AXI_HP2_ID_WIDTH) S_AXI_HP2_RID();
    method Bit#(1) S_AXI_HP2_RLAST();
    method Action S_AXI_HP2_RREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP2_RRESP();
    method Bit#(1) S_AXI_HP2_RVALID();
    method Bit#(6) S_AXI_HP2_WACOUNT();
    method Bit#(8) S_AXI_HP2_WCOUNT();
    method Action S_AXI_HP2_WDATA(Bit#(C_S_AXI_HP2_DATA_WIDTH) v);
    method Action S_AXI_HP2_WID(Bit#(C_S_AXI_HP2_ID_WIDTH) v);
    method Action S_AXI_HP2_WLAST(Bit#(1) v);
    method Bit#(1) S_AXI_HP2_WREADY();
    method Action S_AXI_HP2_WRISSUECAP1_EN(Bit#(1) v);
    method Action S_AXI_HP2_WSTRB(Bit#(C_S_AXI_HP2_DATA_WIDTH) v);
    method Action S_AXI_HP2_WVALID(Bit#(1) v);
    method Action S_AXI_HP3_ACLK(Bit#(1) v);
    method Action S_AXI_HP3_ARADDR(Bit#(32) v);
    method Action S_AXI_HP3_ARBURST(Bit#(2) v);
    method Action S_AXI_HP3_ARCACHE(Bit#(4) v);
    method Bit#(1) S_AXI_HP3_ARESETN();
    method Action S_AXI_HP3_ARID(Bit#(C_S_AXI_HP3_ID_WIDTH) v);
    method Action S_AXI_HP3_ARLEN(Bit#(4) v);
    method Action S_AXI_HP3_ARLOCK(Bit#(2) v);
    method Action S_AXI_HP3_ARPROT(Bit#(3) v);
    method Action S_AXI_HP3_ARQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP3_ARREADY();
    method Action S_AXI_HP3_ARSIZE(Bit#(3) v);
    method Action S_AXI_HP3_ARVALID(Bit#(1) v);
    method Action S_AXI_HP3_AWADDR(Bit#(32) v);
    method Action S_AXI_HP3_AWBURST(Bit#(2) v);
    method Action S_AXI_HP3_AWCACHE(Bit#(4) v);
    method Action S_AXI_HP3_AWID(Bit#(C_S_AXI_HP3_ID_WIDTH) v);
    method Action S_AXI_HP3_AWLEN(Bit#(4) v);
    method Action S_AXI_HP3_AWLOCK(Bit#(2) v);
    method Action S_AXI_HP3_AWPROT(Bit#(3) v);
    method Action S_AXI_HP3_AWQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP3_AWREADY();
    method Action S_AXI_HP3_AWSIZE(Bit#(3) v);
    method Action S_AXI_HP3_AWVALID(Bit#(1) v);
    method Bit#(C_S_AXI_HP3_ID_WIDTH) S_AXI_HP3_BID();
    method Action S_AXI_HP3_BREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP3_BRESP();
    method Bit#(1) S_AXI_HP3_BVALID();
    method Bit#(3) S_AXI_HP3_RACOUNT();
    method Bit#(8) S_AXI_HP3_RCOUNT();
    method Bit#(C_S_AXI_HP3_DATA_WIDTH) S_AXI_HP3_RDATA();
    method Action S_AXI_HP3_RDISSUECAP1_EN(Bit#(1) v);
    method Bit#(C_S_AXI_HP3_ID_WIDTH) S_AXI_HP3_RID();
    method Bit#(1) S_AXI_HP3_RLAST();
    method Action S_AXI_HP3_RREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP3_RRESP();
    method Bit#(1) S_AXI_HP3_RVALID();
    method Bit#(6) S_AXI_HP3_WACOUNT();
    method Bit#(8) S_AXI_HP3_WCOUNT();
    method Action S_AXI_HP3_WDATA(Bit#(C_S_AXI_HP3_DATA_WIDTH) v);
    method Action S_AXI_HP3_WID(Bit#(C_S_AXI_HP3_ID_WIDTH) v);
    method Action S_AXI_HP3_WLAST(Bit#(1) v);
    method Bit#(1) S_AXI_HP3_WREADY();
    method Action S_AXI_HP3_WRISSUECAP1_EN(Bit#(1) v);
    method Action S_AXI_HP3_WSTRB(Bit#(C_S_AXI_HP3_DATA_WIDTH/8) v);
    method Action S_AXI_HP3_WVALID(Bit#(1) v);
    method Action TRACE_CLK(Bit#(1) v);
    method Bit#(1) TRACE_CTL();
    method Bit#(32) TRACE_DATA();
    method Action TTC0_CLK0_IN(Bit#(1) v);
    method Action TTC0_CLK1_IN(Bit#(1) v);
    method Action TTC0_CLK2_IN(Bit#(1) v);
    method Bit#(1) TTC0_WAVE0_OUT();
    method Bit#(1) TTC0_WAVE1_OUT();
    method Bit#(1) TTC0_WAVE2_OUT();
    method Action TTC1_CLK0_IN(Bit#(1) v);
    method Action TTC1_CLK1_IN(Bit#(1) v);
    method Action TTC1_CLK2_IN(Bit#(1) v);
    method Bit#(1) TTC1_WAVE0_OUT();
    method Bit#(1) TTC1_WAVE1_OUT();
    method Bit#(1) TTC1_WAVE2_OUT();
    method Action UART0_CTSN(Bit#(1) v);
    method Action UART0_DCDN(Bit#(1) v);
    method Action UART0_DSRN(Bit#(1) v);
    method Bit#(1) UART0_DTRN();
    method Action UART0_RIN(Bit#(1) v);
    method Bit#(1) UART0_RTSN();
    method Action UART0_RX(Bit#(1) v);
    method Bit#(1) UART0_TX();
    method Action UART1_CTSN(Bit#(1) v);
    method Action UART1_DCDN(Bit#(1) v);
    method Action UART1_DSRN(Bit#(1) v);
    method Bit#(1) UART1_DTRN();
    method Action UART1_RIN(Bit#(1) v);
    method Bit#(1) UART1_RTSN();
    method Action UART1_RX(Bit#(1) v);
    method Bit#(1) UART1_TX();
    method Bit#(2) USB0_PORT_INDCTL();
    method Action USB0_VBUS_PWRFAULT(Bit#(1) v);
    method Bit#(1) USB0_VBUS_PWRSELECT();
    method Bit#(2) USB1_PORT_INDCTL();
    method Action USB1_VBUS_PWRFAULT(Bit#(1) v);
    method Bit#(1) USB1_VBUS_PWRSELECT();
    method Action WDT_CLK_IN(Bit#(1) v);
    method Bit#(1) WDT_RST_OUT();
endinterface

import "BVI" processing_system7 =
module mkPS7(Ps7);
   default_clock clk(C);
   no_reset;
    method Action   (Bit#(1) v); //_clock serdes ()= serdes_clock;

//    parameter USE_TRACE_DATA_EDGE_DETECTOR = 0;
//    parameter C_DM_WIDTH = 0;
//    parameter C_DQS_WIDTH = 0;
//    parameter C_DQ_WIDTH = 0;
//    parameter C_EMIO_GPIO_WIDTH = 0;
//    parameter C_EN_EMIO_ENET0 = 0;
//    parameter C_EN_EMIO_ENET1 = 0;
//    parameter C_EN_EMIO_TRACE = 0;
//    parameter C_FCLK_CLK0_BUF = 0;
//    parameter C_FCLK_CLK1_BUF = 0;
//    parameter C_FCLK_CLK2_BUF = 0;
//    parameter C_FCLK_CLK3_BUF = 0;
//    parameter C_INCLUDE_ACP_TRANS_CHECK = 0;
//    parameter C_INCLUDE_TRACE_BUFFER = 0;
//    parameter C_MIO_PRIMITIVE = 0;
//    parameter C_M_AXI_GP0_ENABLE_STATIC_REMAP = 0;
//    parameter C_M_AXI_GP0_ID_WIDTH = 0;
//    parameter C_M_AXI_GP0_THREAD_ID_WIDTH = 0;
//    parameter C_M_AXI_GP1_ENABLE_STATIC_REMAP = 0;
//    parameter C_M_AXI_GP1_ID_WIDTH = 0;
//    parameter C_M_AXI_GP1_THREAD_ID_WIDTH = 0;
    parameter C_NUM_F2P_INTR_INPUTS = 16;
//    parameter C_PACKAGE_NAME = 0;
//    parameter C_PS7_SI_REV = 0;
//    parameter C_S_AXI_ACP_ARUSER_VAL = 0;
//    parameter C_S_AXI_ACP_AWUSER_VAL = 0;
//    parameter C_S_AXI_ACP_ID_WIDTH = 0;
//    parameter C_S_AXI_GP0_ID_WIDTH = 0;
//    parameter C_S_AXI_GP1_ID_WIDTH = 0;
//    parameter C_S_AXI_HP0_DATA_WIDTH = 0;
//    parameter C_S_AXI_HP0_ID_WIDTH = 0;
//    parameter C_S_AXI_HP1_DATA_WIDTH = 0;
//    parameter C_S_AXI_HP1_ID_WIDTH = 0;
//    parameter C_S_AXI_HP2_DATA_WIDTH = 0;
//    parameter C_S_AXI_HP2_ID_WIDTH = 0;
//    parameter C_S_AXI_HP3_DATA_WIDTH = 0;
//    parameter C_S_AXI_HP3_ID_WIDTH = 0;
//    parameter C_TRACE_BUFFER_CLOCK_DELAY = 0;
//    parameter C_TRACE_BUFFER_FIFO_SIZE = 0;
//    parameter C_USE_DEFAULT_ACP_USER_VAL = 0;

   method CNTVALUEOUT cntvalueout();
   method cinvctrl(CINVCTRL) enable((*inhigh*) en0);
    method Action CAN0_PHY_RX(Bit#(1) v);
    method Bit#(1) CAN0_PHY_TX();
    method Action CAN1_PHY_RX(Bit#(1) v);
    method Bit#(1) CAN1_PHY_TX();
    method Action Core0_nFIQ(Bit#(1) v);
    method Action Core0_nIRQ(Bit#(1) v);
    method Action Core1_nFIQ(Bit#(1) v);
    method Action Core1_nIRQ(Bit#(1) v);
    method Action DDR_ARB(Bit#(4) v);
    method Bit#(15) DDR_Addr();
    method Bit#(3) DDR_BankAddr();
    method Bit#(1) DDR_CAS_n();
    method Bit#(1) DDR_CKE();
    method Bit#(1) DDR_CS_n();
    method Bit#(1) DDR_Clk();
    method Bit#(1) DDR_Clk_n();
    method Bit#(C_DM_WIDTH) DDR_DM();
    method Bit#(C_DQ_WIDTH) DDR_DQ();
    method Bit#(C_DQS_WIDTH) DDR_DQS();
    method Bit#(C_DQS_WIDTH) DDR_DQS_n();
    method Bit#(1) DDR_DRSTB();
    method Bit#(1) DDR_ODT();
    method Bit#(1) DDR_RAS_n();
    method Bit#(1) DDR_VRN();
    method Bit#(1) DDR_VRP();
    method Bit#(1) DDR_WEB();
    method Action DMA0_ACLK(Bit#(1) v);
    method Action DMA0_DAREADY(Bit#(1) v);
    method Bit#(2) DMA0_DATYPE();
    method Bit#(1) DMA0_DAVALID();
    method Action DMA0_DRLAST(Bit#(1) v);
    method Bit#(1) DMA0_DRREADY();
    method Action DMA0_DRTYPE(Bit#(2) v);
    method Action DMA0_DRVALID(Bit#(1) v);
    method Bit#(1) DMA0_RSTN();
    method Action DMA1_ACLK(Bit#(1) v);
    method Action DMA1_DAREADY(Bit#(1) v);
    method Bit#(2) DMA1_DATYPE();
    method Bit#(1) DMA1_DAVALID();
    method Action DMA1_DRLAST(Bit#(1) v);
    method Bit#(1) DMA1_DRREADY();
    method Action DMA1_DRTYPE(Bit#(2) v);
    method Action DMA1_DRVALID(Bit#(1) v);
    method Bit#(1) DMA1_RSTN();
    method Action DMA2_ACLK(Bit#(1) v);
    method Action DMA2_DAREADY(Bit#(1) v);
    method Bit#(2) DMA2_DATYPE();
    method Bit#(1) DMA2_DAVALID();
    method Action DMA2_DRLAST(Bit#(1) v);
    method Bit#(1) DMA2_DRREADY();
    method Action DMA2_DRTYPE(Bit#(2) v);
    method Action DMA2_DRVALID(Bit#(1) v);
    method Bit#(1) DMA2_RSTN();
    method Action DMA3_ACLK(Bit#(1) v);
    method Action DMA3_DAREADY(Bit#(1) v);
    method Bit#(2) DMA3_DATYPE();
    method Bit#(1) DMA3_DAVALID();
    method Action DMA3_DRLAST(Bit#(1) v);
    method Bit#(1) DMA3_DRREADY();
    method Action DMA3_DRTYPE(Bit#(2) v);
    method Action DMA3_DRVALID(Bit#(1) v);
    method Bit#(1) DMA3_RSTN();
    method Action ENET0_EXT_INTIN(Bit#(1) v);
    method Action ENET0_GMII_COL(Bit#(1) v);
    method Action ENET0_GMII_CRS(Bit#(1) v);
    method Action ENET0_GMII_RXD(Bit#(8) v);
    method Action ENET0_GMII_RX_CLK(Bit#(1) v);
    method Action ENET0_GMII_RX_DV(Bit#(1) v);
    method Action ENET0_GMII_RX_ER(Bit#(1) v);
    method Bit#(8) ENET0_GMII_TXD();
    method Action ENET0_GMII_TX_CLK(Bit#(1) v);
    method Bit#(1) ENET0_GMII_TX_EN();
    method Bit#(1) ENET0_GMII_TX_ER();
    method Action ENET0_MDIO_I(Bit#(1) v);
    method Bit#(1) ENET0_MDIO_MDC();
    method Bit#(1) ENET0_MDIO_O();
    method Bit#(1) ENET0_MDIO_T();
    method Bit#(1) ENET0_PTP_DELAY_REQ_RX();
    method Bit#(1) ENET0_PTP_DELAY_REQ_TX();
    method Bit#(1) ENET0_PTP_PDELAY_REQ_RX();
    method Bit#(1) ENET0_PTP_PDELAY_REQ_TX();
    method Bit#(1) ENET0_PTP_PDELAY_RESP_RX();
    method Bit#(1) ENET0_PTP_PDELAY_RESP_TX();
    method Bit#(1) ENET0_PTP_SYNC_FRAME_RX();
    method Bit#(1) ENET0_PTP_SYNC_FRAME_TX();
    method Bit#(1) ENET0_SOF_RX();
    method Bit#(1) ENET0_SOF_TX();
    method Action ENET1_EXT_INTIN(Bit#(1) v);
    method Action ENET1_GMII_COL(Bit#(1) v);
    method Action ENET1_GMII_CRS(Bit#(1) v);
    method Action ENET1_GMII_RXD(Bit#(8) v);
    method Action ENET1_GMII_RX_CLK(Bit#(1) v);
    method Action ENET1_GMII_RX_DV(Bit#(1) v);
    method Action ENET1_GMII_RX_ER(Bit#(1) v);
    method Bit#(8) ENET1_GMII_TXD();
    method Action ENET1_GMII_TX_CLK(Bit#(1) v);
    method Bit#(1) ENET1_GMII_TX_EN();
    method Bit#(1) ENET1_GMII_TX_ER();
    method Action ENET1_MDIO_I(Bit#(1) v);
    method Bit#(1) ENET1_MDIO_MDC();
    method Bit#(1) ENET1_MDIO_O();
    method Bit#(1) ENET1_MDIO_T();
    method Bit#(1) ENET1_PTP_DELAY_REQ_RX();
    method Bit#(1) ENET1_PTP_DELAY_REQ_TX();
    method Bit#(1) ENET1_PTP_PDELAY_REQ_RX();
    method Bit#(1) ENET1_PTP_PDELAY_REQ_TX();
    method Bit#(1) ENET1_PTP_PDELAY_RESP_RX();
    method Bit#(1) ENET1_PTP_PDELAY_RESP_TX();
    method Bit#(1) ENET1_PTP_SYNC_FRAME_RX();
    method Bit#(1) ENET1_PTP_SYNC_FRAME_TX();
    method Bit#(1) ENET1_SOF_RX();
    method Bit#(1) ENET1_SOF_TX();
    method Action EVENT_EVENTI(Bit#(1) v);
    method Bit#(1) EVENT_EVENTO();
    method Bit#(2) EVENT_STANDBYWFE();
    method Bit#(2) EVENT_STANDBYWFI();
    method Bit#(1) FCLK_CLK0();
    method Bit#(1) FCLK_CLK1();
    method Bit#(1) FCLK_CLK2();
    method Bit#(1) FCLK_CLK3();
    method Action FCLK_CLKTRIG0_N(Bit#(1) v);
    method Action FCLK_CLKTRIG1_N(Bit#(1) v);
    method Action FCLK_CLKTRIG2_N(Bit#(1) v);
    method Action FCLK_CLKTRIG3_N(Bit#(1) v);
    method Bit#(1) FCLK_RESET0_N();
    method Bit#(1) FCLK_RESET1_N();
    method Bit#(1) FCLK_RESET2_N();
    method Bit#(1) FCLK_RESET3_N();
    method Action FPGA_IDLE_N(Bit#(1) v);
    method Action FTMD_TRACEIN_ATID(Bit#(4) v);
    method Action FTMD_TRACEIN_CLK(Bit#(1) v);
    method Action FTMD_TRACEIN_DATA(Bit#(32) v);
    method Action FTMD_TRACEIN_VALID(Bit#(1) v);
    method Action FTMT_F2P_DEBUG(Bit#(32) v);
    method Action FTMT_F2P_TRIG(Bit#(4) v);
    method Bit#(4) FTMT_F2P_TRIGACK();
    method Bit#(32) FTMT_P2F_DEBUG();
    method Bit#(4) FTMT_P2F_TRIG();
    method Action FTMT_P2F_TRIGACK(Bit#(4) v);
    method Action GPIO_I(Bit#(C_EMIO_GPIO_WIDTH) v);
    method Bit#(C_EMIO_GPIO_WIDTH) GPIO_O();
    method Bit#(C_EMIO_GPIO_WIDTH) GPIO_T();
    method Action I2C0_SCL_I(Bit#(1) v);
    method Bit#(1) I2C0_SCL_O();
    method Bit#(1) I2C0_SCL_T();
    method Action I2C0_SDA_I(Bit#(1) v);
    method Bit#(1) I2C0_SDA_O();
    method Bit#(1) I2C0_SDA_T();
    method Action I2C1_SCL_I(Bit#(1) v);
    method Bit#(1) I2C1_SCL_O();
    method Bit#(1) I2C1_SCL_T();
    method Action I2C1_SDA_I(Bit#(1) v);
    method Bit#(1) I2C1_SDA_O();
    method Bit#(1) I2C1_SDA_T();
    method Action IRQ_F2P(Bit#(16) v);
    method Bit#(1) IRQ_P2F_CAN0();
    method Bit#(1) IRQ_P2F_CAN1();
    method Bit#(1) IRQ_P2F_CTI();
    method Bit#(1) IRQ_P2F_DMAC0();
    method Bit#(1) IRQ_P2F_DMAC1();
    method Bit#(1) IRQ_P2F_DMAC2();
    method Bit#(1) IRQ_P2F_DMAC3();
    method Bit#(1) IRQ_P2F_DMAC4();
    method Bit#(1) IRQ_P2F_DMAC5();
    method Bit#(1) IRQ_P2F_DMAC6();
    method Bit#(1) IRQ_P2F_DMAC7();
    method Bit#(1) IRQ_P2F_DMAC_ABORT();
    method Bit#(1) IRQ_P2F_ENET0();
    method Bit#(1) IRQ_P2F_ENET1();
    method Bit#(1) IRQ_P2F_ENET_WAKE0();
    method Bit#(1) IRQ_P2F_ENET_WAKE1();
    method Bit#(1) IRQ_P2F_GPIO();
    method Bit#(1) IRQ_P2F_I2C0();
    method Bit#(1) IRQ_P2F_I2C1();
    method Bit#(1) IRQ_P2F_QSPI();
    method Bit#(1) IRQ_P2F_SDIO0();
    method Bit#(1) IRQ_P2F_SDIO1();
    method Bit#(1) IRQ_P2F_SMC();
    method Bit#(1) IRQ_P2F_SPI0();
    method Bit#(1) IRQ_P2F_SPI1();
    method Bit#(1) IRQ_P2F_UART0();
    method Bit#(1) IRQ_P2F_UART1();
    method Bit#(1) IRQ_P2F_USB0();
    method Bit#(1) IRQ_P2F_USB1();
    method Bit#(C_MIO_PRIMITIVE) MIO();
    method Action M_AXI_GP0_ACLK(Bit#(1) v);
    method Bit#(32) M_AXI_GP0_ARADDR();
    method Bit#(2) M_AXI_GP0_ARBURST();
    method Bit#(4) M_AXI_GP0_ARCACHE();
    method Bit#(1) M_AXI_GP0_ARESETN();
    method Bit#(C_M_AXI_GP0_THREAD_ID_WIDTH) M_AXI_GP0_ARID();
    method Bit#(4) M_AXI_GP0_ARLEN();
    method Bit#(2) M_AXI_GP0_ARLOCK();
    method Bit#(3) M_AXI_GP0_ARPROT();
    method Bit#(4) M_AXI_GP0_ARQOS();
    method Action M_AXI_GP0_ARREADY(Bit#(1) v);
    method Bit#(3) M_AXI_GP0_ARSIZE();
    method Bit#(1) M_AXI_GP0_ARVALID();
    method Bit#(32) M_AXI_GP0_AWADDR();
    method Bit#(2) M_AXI_GP0_AWBURST();
    method Bit#(4) M_AXI_GP0_AWCACHE();
    method Bit#(C_M_AXI_GP0_THREAD_ID_WIDTH) M_AXI_GP0_AWID();
    method Bit#(4) M_AXI_GP0_AWLEN();
    method Bit#(2) M_AXI_GP0_AWLOCK();
    method Bit#(3) M_AXI_GP0_AWPROT();
    method Bit#(4) M_AXI_GP0_AWQOS();
    method Action M_AXI_GP0_AWREADY(Bit#(1) v);
    method Bit#(3) M_AXI_GP0_AWSIZE();
    method Bit#(1) M_AXI_GP0_AWVALID();
    method Action M_AXI_GP0_BID(Bit#(C_M_AXI_GP0_THREAD_ID_WIDTH) v);
    method Bit#(1) M_AXI_GP0_BREADY();
    method Action M_AXI_GP0_BRESP(Bit#(2) v);
    method Action M_AXI_GP0_BVALID(Bit#(1) v);
    method Action M_AXI_GP0_RDATA(Bit#(32) v);
    method Action M_AXI_GP0_RID(Bit#(C_M_AXI_GP0_THREAD_ID_WIDTH) v);
    method Action M_AXI_GP0_RLAST(Bit#(1) v);
    method Bit#(1) M_AXI_GP0_RREADY();
    method Action M_AXI_GP0_RRESP(Bit#(2) v);
    method Action M_AXI_GP0_RVALID(Bit#(1) v);
    method Bit#(32) M_AXI_GP0_WDATA();
    method Bit#(C_M_AXI_GP0_THREAD_ID_WIDTH) M_AXI_GP0_WID();
    method Bit#(1) M_AXI_GP0_WLAST();
    method Action M_AXI_GP0_WREADY(Bit#(1) v);
    method Bit#(4) M_AXI_GP0_WSTRB();
    method Bit#(1) M_AXI_GP0_WVALID();
    method Action M_AXI_GP1_ACLK(Bit#(1) v);
    method Bit#(32) M_AXI_GP1_ARADDR();
    method Bit#(2) M_AXI_GP1_ARBURST();
    method Bit#(4) M_AXI_GP1_ARCACHE();
    method Bit#(1) M_AXI_GP1_ARESETN();
    method Bit#(C_M_AXI_GP1_THREAD_ID_WIDTH) M_AXI_GP1_ARID();
    method Bit#(4) M_AXI_GP1_ARLEN();
    method Bit#(2) M_AXI_GP1_ARLOCK();
    method Bit#(3) M_AXI_GP1_ARPROT();
    method Bit#(4) M_AXI_GP1_ARQOS();
    method Action M_AXI_GP1_ARREADY(Bit#(1) v);
    method Bit#(3) M_AXI_GP1_ARSIZE();
    method Bit#(1) M_AXI_GP1_ARVALID();
    method Bit#(32) M_AXI_GP1_AWADDR();
    method Bit#(2) M_AXI_GP1_AWBURST();
    method Bit#(4) M_AXI_GP1_AWCACHE();
    method Bit#(C_M_AXI_GP1_THREAD_ID_WIDTH) M_AXI_GP1_AWID();
    method Bit#(4) M_AXI_GP1_AWLEN();
    method Bit#(2) M_AXI_GP1_AWLOCK();
    method Bit#(3) M_AXI_GP1_AWPROT();
    method Bit#(4) M_AXI_GP1_AWQOS();
    method Action M_AXI_GP1_AWREADY(Bit#(1) v);
    method Bit#(3) M_AXI_GP1_AWSIZE();
    method Bit#(1) M_AXI_GP1_AWVALID();
    method Action M_AXI_GP1_BID(Bit#(C_M_AXI_GP1_THREAD_ID_WIDTH) v);
    method Bit#(1) M_AXI_GP1_BREADY();
    method Action M_AXI_GP2_BRESP(Bit#(1) v);
    method Action M_AXI_GP1_BVALID(Bit#(1) v);
    method Action M_AXI_GP1_RDATA(Bit#(32) v);
    method Action M_AXI_GP1_RID(Bit#(C_M_AXI_GP1_THREAD_ID_WIDTH) v);
    method Action M_AXI_GP1_RLAST(Bit#(1) v);
    method Bit#(1) M_AXI_GP1_RREADY();
    method Action M_AXI_GP2_RRESP(Bit#(1) v);
    method Action M_AXI_GP1_RVALID(Bit#(1) v);
    method Bit#(32) M_AXI_GP1_WDATA();
    method Bit#(C_M_AXI_GP1_THREAD_ID_WIDTH) M_AXI_GP1_WID();
    method Bit#(1) M_AXI_GP1_WLAST();
    method Action M_AXI_GP1_WREADY(Bit#(1) v);
    method Bit#(4) M_AXI_GP1_WSTRB();
    method Bit#(1) M_AXI_GP1_WVALID();
    method Action PJTAG_TCK(Bit#(1) v);
    method Action PJTAG_TD_I(Bit#(1) v);
    method Bit#(1) PJTAG_TD_O();
    method Bit#(1) PJTAG_TD_T();
    method Action PJTAG_TMS(Bit#(1) v);
    method Action PS_CLK(Bit#(1) v);
    method Action PS_PORB(Bit#(1) v);
    method Action PS_SRSTB(Bit#(1) v);
    method Bit#(1) SDIO0_BUSPOW();
    method Bit#(3) SDIO0_BUSVOLT();
    method Action SDIO0_CDN(Bit#(1) v);
    method Bit#(1) SDIO0_CLK();
    method Action SDIO0_CLK_FB(Bit#(1) v);
    method Action SDIO0_CMD_I(Bit#(1) v);
    method Bit#(1) SDIO0_CMD_O();
    method Bit#(1) SDIO0_CMD_T();
    method Action SDIO0_DATA_I(Bit#(4) v);
    method Bit#(4) SDIO0_DATA_O();
    method Bit#(4) SDIO0_DATA_T();
    method Bit#(1) SDIO0_LED();
    method Action SDIO0_WP(Bit#(1) v);
    method Bit#(1) SDIO1_BUSPOW();
    method Bit#(3) SDIO1_BUSVOLT();
    method Action SDIO1_CDN(Bit#(1) v);
    method Bit#(1) SDIO1_CLK();
    method Action SDIO1_CLK_FB(Bit#(1) v);
    method Action SDIO1_CMD_I(Bit#(1) v);
    method Bit#(1) SDIO1_CMD_O();
    method Bit#(1) SDIO1_CMD_T();
    method Action SDIO1_DATA_I(Bit#(4) v);
    method Bit#(4) SDIO1_DATA_O();
    method Bit#(4) SDIO1_DATA_T();
    method Bit#(1) SDIO1_LED();
    method Action SDIO1_WP(Bit#(1) v);
    method Action SPI0_MISO_I(Bit#(1) v);
    method Bit#(1) SPI0_MISO_O();
    method Bit#(1) SPI0_MISO_T();
    method Action SPI0_MOSI_I(Bit#(1) v);
    method Bit#(1) SPI0_MOSI_O();
    method Bit#(1) SPI0_MOSI_T();
    method Action SPI0_SCLK_I(Bit#(1) v);
    method Bit#(1) SPI0_SCLK_O();
    method Bit#(1) SPI0_SCLK_T();
    method Bit#(1) SPI0_SS1_O();
    method Bit#(1) SPI0_SS2_O();
    method Action SPI0_SS_I(Bit#(1) v);
    method Bit#(1) SPI0_SS_O();
    method Bit#(1) SPI0_SS_T();
    method Action SPI1_MISO_I(Bit#(1) v);
    method Bit#(1) SPI1_MISO_O();
    method Bit#(1) SPI1_MISO_T();
    method Action SPI1_MOSI_I(Bit#(1) v);
    method Bit#(1) SPI1_MOSI_O();
    method Bit#(1) SPI1_MOSI_T();
    method Action SPI1_SCLK_I(Bit#(1) v);
    method Bit#(1) SPI1_SCLK_O();
    method Bit#(1) SPI1_SCLK_T();
    method Bit#(1) SPI1_SS1_O();
    method Bit#(1) SPI1_SS2_O();
    method Action SPI1_SS_I(Bit#(1) v);
    method Bit#(1) SPI1_SS_O();
    method Bit#(1) SPI1_SS_T();
    method Action SRAM_INTIN(Bit#(1) v);
    method Action S_AXI_ACP_ACLK(Bit#(1) v);
    method Action S_AXI_ACP_ARADDR(Bit#(32) v);
    method Action S_AXI_ACP_ARBURST(Bit#(2) v);
    method Action S_AXI_ACP_ARCACHE(Bit#(4) v);
    method Bit#(1) S_AXI_ACP_ARESETN();
    method Action S_AXI_ACP_ARID(Bit#(C_S_AXI_ACP_ID_WIDTH) v);
    method Action S_AXI_ACP_ARLEN(Bit#(4) v);
    method Action S_AXI_ACP_ARLOCK(Bit#(2) v);
    method Action S_AXI_ACP_ARPROT(Bit#(3) v);
    method Action S_AXI_ACP_ARQOS(Bit#(4) v);
    method Bit#(1) S_AXI_ACP_ARREADY();
    method Action S_AXI_ACP_ARSIZE(Bit#(3) v);
    method Action S_AXI_ACP_ARUSER(Bit#(5) v);
    method Action S_AXI_ACP_ARVALID(Bit#(1) v);
    method Action S_AXI_ACP_AWADDR(Bit#(32) v);
    method Action S_AXI_ACP_AWBURST(Bit#(2) v);
    method Action S_AXI_ACP_AWCACHE(Bit#(4) v);
    method Action S_AXI_ACP_AWID(Bit#(C_S_AXI_ACP_ID_WIDTH) v);
    method Action S_AXI_ACP_AWLEN(Bit#(4) v);
    method Action S_AXI_ACP_AWLOCK(Bit#(2) v);
    method Action S_AXI_ACP_AWPROT(Bit#(3) v);
    method Action S_AXI_ACP_AWQOS(Bit#(4) v);
    method Bit#(1) S_AXI_ACP_AWREADY();
    method Action S_AXI_ACP_AWSIZE(Bit#(3) v);
    method Action S_AXI_ACP_AWUSER(Bit#(5) v);
    method Action S_AXI_ACP_AWVALID(Bit#(1) v);
    method Bit#(C_S_AXI_ACP_ID_WIDTH) S_AXI_ACP_BID();
    method Action S_AXI_ACP_BREADY(Bit#(1) v);
    method Bit#(2) S_AXI_ACP_BRESP();
    method Bit#(1) S_AXI_ACP_BVALID();
    method Bit#(64) S_AXI_ACP_RDATA();
    method Bit#(C_S_AXI_ACP_ID_WIDTH) S_AXI_ACP_RID();
    method Bit#(1) S_AXI_ACP_RLAST();
    method Action S_AXI_ACP_RREADY(Bit#(1) v);
    method Bit#(2) S_AXI_ACP_RRESP();
    method Bit#(1) S_AXI_ACP_RVALID();
    method Action S_AXI_ACP_WDATA(Bit#(64) v);
    method Action S_AXI_ACP_WID(Bit#(C_S_AXI_ACP_ID_WIDTH) v);
    method Action S_AXI_ACP_WLAST(Bit#(1) v);
    method Bit#(1) S_AXI_ACP_WREADY();
    method Action S_AXI_ACP_WSTRB(Bit#(8) v);
    method Action S_AXI_ACP_WVALID(Bit#(1) v);
    method Action S_AXI_GP0_ACLK(Bit#(1) v);
    method Action S_AXI_GP0_ARADDR(Bit#(32) v);
    method Action S_AXI_GP0_ARBURST(Bit#(2) v);
    method Action S_AXI_GP0_ARCACHE(Bit#(4) v);
    method Bit#(1) S_AXI_GP0_ARESETN();
    method Action S_AXI_GP0_ARID(Bit#(C_S_AXI_GP0_ID_WIDTH) v);
    method Action S_AXI_GP0_ARLEN(Bit#(4) v);
    method Action S_AXI_GP0_ARLOCK(Bit#(2) v);
    method Action S_AXI_GP0_ARPROT(Bit#(3) v);
    method Action S_AXI_GP0_ARQOS(Bit#(4) v);
    method Bit#(1) S_AXI_GP0_ARREADY();
    method Action S_AXI_GP0_ARSIZE(Bit#(3) v);
    method Action S_AXI_GP0_ARVALID(Bit#(1) v);
    method Action S_AXI_GP0_AWADDR(Bit#(32) v);
    method Action S_AXI_GP0_AWBURST(Bit#(2) v);
    method Action S_AXI_GP0_AWCACHE(Bit#(4) v);
    method Action S_AXI_GP0_AWID(Bit#(C_S_AXI_GP0_ID_WIDTH) v);
    method Action S_AXI_GP0_AWLEN(Bit#(4) v);
    method Action S_AXI_GP0_AWLOCK(Bit#(2) v);
    method Action S_AXI_GP0_AWPROT(Bit#(3) v);
    method Action S_AXI_GP0_AWQOS(Bit#(4) v);
    method Bit#(1) S_AXI_GP0_AWREADY();
    method Action S_AXI_GP0_AWSIZE(Bit#(3) v);
    method Action S_AXI_GP0_AWVALID(Bit#(1) v);
    method Bit#(C_S_AXI_GP0_ID_WIDTH) S_AXI_GP0_BID();
    method Action S_AXI_GP0_BREADY(Bit#(1) v);
    method Bit#(2) S_AXI_GP0_BRESP();
    method Bit#(1) S_AXI_GP0_BVALID();
    method Bit#(32) S_AXI_GP0_RDATA();
    method Bit#(C_S_AXI_GP0_ID_WIDTH) S_AXI_GP0_RID();
    method Bit#(1) S_AXI_GP0_RLAST();
    method Action S_AXI_GP0_RREADY(Bit#(1) v);
    method Bit#(2) S_AXI_GP0_RRESP();
    method Bit#(1) S_AXI_GP0_RVALID();
    method Action S_AXI_GP0_WDATA(Bit#(32) v);
    method Action S_AXI_GP0_WID(Bit#(C_S_AXI_GP0_ID_WIDTH) v);
    method Action S_AXI_GP0_WLAST(Bit#(1) v);
    method Bit#(1) S_AXI_GP0_WREADY();
    method Action S_AXI_GP0_WSTRB(Bit#(4) v);
    method Action S_AXI_GP0_WVALID(Bit#(1) v);
    method Action S_AXI_GP1_ACLK(Bit#(1) v);
    method Action S_AXI_GP1_ARADDR(Bit#(32) v);
    method Action S_AXI_GP2_ARBURST(Bit#(1) v);
    method Action S_AXI_GP1_ARCACHE(Bit#(4) v);
    method Bit#(1) S_AXI_GP1_ARESETN();
    method Action S_AXI_GP1_ARID(Bit#(C_S_AXI_GP1_ID_WIDTH) v);
    method Action S_AXI_GP1_ARLEN(Bit#(4) v);
    method Action S_AXI_GP2_ARLOCK(Bit#(1) v);
    method Action S_AXI_GP1_ARPROT(Bit#(3) v);
    method Action S_AXI_GP1_ARQOS(Bit#(4) v);
    method Bit#(1) S_AXI_GP1_ARREADY();
    method Action S_AXI_GP1_ARSIZE(Bit#(3) v);
    method Action S_AXI_GP1_ARVALID(Bit#(1) v);
    method Action S_AXI_GP1_AWADDR(Bit#(32) v);
    method Action S_AXI_GP2_AWBURST(Bit#(1) v);
    method Action S_AXI_GP1_AWCACHE(Bit#(4) v);
    method Action S_AXI_GP1_AWID(Bit#(C_S_AXI_GP1_ID_WIDTH) v);
    method Action S_AXI_GP1_AWLEN(Bit#(4) v);
    method Action S_AXI_GP2_AWLOCK(Bit#(1) v);
    method Action S_AXI_GP1_AWPROT(Bit#(3) v);
    method Action S_AXI_GP1_AWQOS(Bit#(4) v);
    method Bit#(1) S_AXI_GP1_AWREADY();
    method Action S_AXI_GP1_AWSIZE(Bit#(3) v);
    method Action S_AXI_GP1_AWVALID(Bit#(1) v);
    method Bit#(C_S_AXI_GP1_ID_WIDTH) S_AXI_GP1_BID();
    method Action S_AXI_GP1_BREADY(Bit#(1) v);
    method Bit#(2) S_AXI_GP1_BRESP();
    method Bit#(1) S_AXI_GP1_BVALID();
    method Bit#(32) S_AXI_GP1_RDATA();
    method Bit#(C_S_AXI_GP1_ID_WIDTH) S_AXI_GP1_RID();
    method Bit#(1) S_AXI_GP1_RLAST();
    method Action S_AXI_GP1_RREADY(Bit#(1) v);
    method Bit#(2) S_AXI_GP1_RRESP();
    method Bit#(1) S_AXI_GP1_RVALID();
    method Action S_AXI_GP1_WDATA(Bit#(32) v);
    method Action S_AXI_GP1_WID(Bit#(C_S_AXI_GP1_ID_WIDTH) v);
    method Action S_AXI_GP1_WLAST(Bit#(1) v);
    method Bit#(1) S_AXI_GP1_WREADY();
    method Action S_AXI_GP1_WSTRB(Bit#(4) v);
    method Action S_AXI_GP1_WVALID(Bit#(1) v);
    method Action S_AXI_HP0_ACLK(Bit#(1) v);
    method Action S_AXI_HP0_ARADDR(Bit#(32) v);
    method Action S_AXI_HP0_ARBURST(Bit#(2) v);
    method Action S_AXI_HP0_ARCACHE(Bit#(4) v);
    method Bit#(1) S_AXI_HP0_ARESETN();
    method Action S_AXI_HP0_ARID(Bit#(C_S_AXI_HP0_ID_WIDTH) v);
    method Action S_AXI_HP0_ARLEN(Bit#(4) v);
    method Action S_AXI_HP0_ARLOCK(Bit#(2) v);
    method Action S_AXI_HP0_ARPROT(Bit#(3) v);
    method Action S_AXI_HP0_ARQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP0_ARREADY();
    method Action S_AXI_HP0_ARSIZE(Bit#(3) v);
    method Action S_AXI_HP0_ARVALID(Bit#(1) v);
    method Action S_AXI_HP0_AWADDR(Bit#(32) v);
    method Action S_AXI_HP0_AWBURST(Bit#(2) v);
    method Action S_AXI_HP0_AWCACHE(Bit#(4) v);
    method Action S_AXI_HP0_AWID(Bit#(C_S_AXI_HP0_ID_WIDTH) v);
    method Action S_AXI_HP0_AWLEN(Bit#(4) v);
    method Action S_AXI_HP0_AWLOCK(Bit#(2) v);
    method Action S_AXI_HP0_AWPROT(Bit#(3) v);
    method Action S_AXI_HP0_AWQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP0_AWREADY();
    method Action S_AXI_HP0_AWSIZE(Bit#(3) v);
    method Action S_AXI_HP0_AWVALID(Bit#(1) v);
    method Bit#(C_S_AXI_HP0_ID_WIDTH) S_AXI_HP0_BID();
    method Action S_AXI_HP0_BREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP0_BRESP();
    method Bit#(1) S_AXI_HP0_BVALID();
    method Bit#(3) S_AXI_HP0_RACOUNT();
    method Bit#(8) S_AXI_HP0_RCOUNT();
    method Bit#(C_S_AXI_HP0_DATA_WIDTH) S_AXI_HP0_RDATA();
    method Action S_AXI_HP0_RDISSUECAP1_EN(Bit#(1) v);
    method Bit#(C_S_AXI_HP0_ID_WIDTH) S_AXI_HP0_RID();
    method Bit#(1) S_AXI_HP0_RLAST();
    method Action S_AXI_HP0_RREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP0_RRESP();
    method Bit#(1) S_AXI_HP0_RVALID();
    method Bit#(6) S_AXI_HP0_WACOUNT();
    method Bit#(8) S_AXI_HP0_WCOUNT();
    method Action S_AXI_HP0_WDATA(Bit#(C_S_AXI_HP0_DATA_WIDTH) v);
    method Action S_AXI_HP0_WID(Bit#(C_S_AXI_HP0_ID_WIDTH) v);
    method Action S_AXI_HP0_WLAST(Bit#(1) v);
    method Bit#(1) S_AXI_HP0_WREADY();
    method Action S_AXI_HP0_WRISSUECAP1_EN(Bit#(1) v);
    method Action S_AXI_HP0_WSTRB(Bit#(C_S_AXI_HP0_DATA_WIDTH/8) v);
    method Action S_AXI_HP0_WVALID(Bit#(1) v);
    method Action S_AXI_HP1_ACLK(Bit#(1) v);
    method Action S_AXI_HP1_ARADDR(Bit#(32) v);
    method Action S_AXI_HP2_ARBURST(Bit#(1) v);
    method Action S_AXI_HP1_ARCACHE(Bit#(4) v);
    method Bit#(1) S_AXI_HP1_ARESETN();
    method Action S_AXI_HP1_ARID(Bit#(C_S_AXI_HP1_ID_WIDTH) v);
    method Action S_AXI_HP1_ARLEN(Bit#(4) v);
    method Action S_AXI_HP2_ARLOCK(Bit#(1) v);
    method Action S_AXI_HP1_ARPROT(Bit#(3) v);
    method Action S_AXI_HP1_ARQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP1_ARREADY();
    method Action S_AXI_HP1_ARSIZE(Bit#(3) v);
    method Action S_AXI_HP1_ARVALID(Bit#(1) v);
    method Action S_AXI_HP1_AWADDR(Bit#(32) v);
    method Action S_AXI_HP2_AWBURST(Bit#(1) v);
    method Action S_AXI_HP1_AWCACHE(Bit#(4) v);
    method Action S_AXI_HP1_AWID(Bit#(C_S_AXI_HP1_ID_WIDTH) v);
    method Action S_AXI_HP1_AWLEN(Bit#(4) v);
    method Action S_AXI_HP2_AWLOCK(Bit#(1) v);
    method Action S_AXI_HP1_AWPROT(Bit#(3) v);
    method Action S_AXI_HP1_AWQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP1_AWREADY();
    method Action S_AXI_HP1_AWSIZE(Bit#(3) v);
    method Action S_AXI_HP1_AWVALID(Bit#(1) v);
    method Bit#(C_S_AXI_HP1_ID_WIDTH) S_AXI_HP1_BID();
    method Action S_AXI_HP1_BREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP1_BRESP();
    method Bit#(1) S_AXI_HP1_BVALID();
    method Bit#(3) S_AXI_HP1_RACOUNT();
    method Bit#(8) S_AXI_HP1_RCOUNT();
    method Bit#(C_S_AXI_HP1_DATA_WIDTH) S_AXI_HP1_RDATA();
    method Action S_AXI_HP1_RDISSUECAP1_EN(Bit#(1) v);
    method Bit#(C_S_AXI_HP1_ID_WIDTH) S_AXI_HP1_RID();
    method Bit#(1) S_AXI_HP1_RLAST();
    method Action S_AXI_HP1_RREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP1_RRESP();
    method Bit#(1) S_AXI_HP1_RVALID();
    method Bit#(6) S_AXI_HP1_WACOUNT();
    method Bit#(8) S_AXI_HP1_WCOUNT();
    method Action S_AXI_HP1_WDATA(Bit#(C_S_AXI_HP1_DATA_WIDTH) v);
    method Action S_AXI_HP1_WID(Bit#(C_S_AXI_HP1_ID_WIDTH) v);
    method Action S_AXI_HP1_WLAST(Bit#(1) v);
    method Bit#(1) S_AXI_HP1_WREADY();
    method Action S_AXI_HP1_WRISSUECAP1_EN(Bit#(1) v);
    method Action S_AXI_HP1_WSTRB(Bit#(C_S_AXI_HP1_DATA_WIDTH) v);
    method Action S_AXI_HP1_WVALID(Bit#(1) v);
    method Action S_AXI_HP2_ACLK(Bit#(1) v);
    method Action S_AXI_HP2_ARADDR(Bit#(32) v);
    method Action S_AXI_HP2_ARBURST(Bit#(2) v);
    method Action S_AXI_HP2_ARCACHE(Bit#(4) v);
    method Bit#(1) S_AXI_HP2_ARESETN();
    method Action S_AXI_HP2_ARID(Bit#(C_S_AXI_HP2_ID_WIDTH) v);
    method Action S_AXI_HP2_ARLEN(Bit#(4) v);
    method Action S_AXI_HP2_ARLOCK(Bit#(2) v);
    method Action S_AXI_HP2_ARPROT(Bit#(3) v);
    method Action S_AXI_HP2_ARQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP2_ARREADY();
    method Action S_AXI_HP2_ARSIZE(Bit#(3) v);
    method Action S_AXI_HP2_ARVALID(Bit#(1) v);
    method Action S_AXI_HP2_AWADDR(Bit#(32) v);
    method Action S_AXI_HP2_AWBURST(Bit#(2) v);
    method Action S_AXI_HP2_AWCACHE(Bit#(4) v);
    method Action S_AXI_HP2_AWID(Bit#(C_S_AXI_HP2_ID_WIDTH) v);
    method Action S_AXI_HP2_AWLEN(Bit#(4) v);
    method Action S_AXI_HP2_AWLOCK(Bit#(2) v);
    method Action S_AXI_HP2_AWPROT(Bit#(3) v);
    method Action S_AXI_HP2_AWQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP2_AWREADY();
    method Action S_AXI_HP2_AWSIZE(Bit#(3) v);
    method Action S_AXI_HP2_AWVALID(Bit#(1) v);
    method Bit#(C_S_AXI_HP2_ID_WIDTH) S_AXI_HP2_BID();
    method Action S_AXI_HP2_BREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP2_BRESP();
    method Bit#(1) S_AXI_HP2_BVALID();
    method Bit#(3) S_AXI_HP2_RACOUNT();
    method Bit#(8) S_AXI_HP2_RCOUNT();
    method Bit#(C_S_AXI_HP2_DATA_WIDTH) S_AXI_HP2_RDATA();
    method Action S_AXI_HP2_RDISSUECAP1_EN(Bit#(1) v);
    method Bit#(C_S_AXI_HP2_ID_WIDTH) S_AXI_HP2_RID();
    method Bit#(1) S_AXI_HP2_RLAST();
    method Action S_AXI_HP2_RREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP2_RRESP();
    method Bit#(1) S_AXI_HP2_RVALID();
    method Bit#(6) S_AXI_HP2_WACOUNT();
    method Bit#(8) S_AXI_HP2_WCOUNT();
    method Action S_AXI_HP2_WDATA(Bit#(C_S_AXI_HP2_DATA_WIDTH) v);
    method Action S_AXI_HP2_WID(Bit#(C_S_AXI_HP2_ID_WIDTH) v);
    method Action S_AXI_HP2_WLAST(Bit#(1) v);
    method Bit#(1) S_AXI_HP2_WREADY();
    method Action S_AXI_HP2_WRISSUECAP1_EN(Bit#(1) v);
    method Action S_AXI_HP2_WSTRB(Bit#(C_S_AXI_HP2_DATA_WIDTH) v);
    method Action S_AXI_HP2_WVALID(Bit#(1) v);
    method Action S_AXI_HP3_ACLK(Bit#(1) v);
    method Action S_AXI_HP3_ARADDR(Bit#(32) v);
    method Action S_AXI_HP3_ARBURST(Bit#(2) v);
    method Action S_AXI_HP3_ARCACHE(Bit#(4) v);
    method Bit#(1) S_AXI_HP3_ARESETN();
    method Action S_AXI_HP3_ARID(Bit#(C_S_AXI_HP3_ID_WIDTH) v);
    method Action S_AXI_HP3_ARLEN(Bit#(4) v);
    method Action S_AXI_HP3_ARLOCK(Bit#(2) v);
    method Action S_AXI_HP3_ARPROT(Bit#(3) v);
    method Action S_AXI_HP3_ARQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP3_ARREADY();
    method Action S_AXI_HP3_ARSIZE(Bit#(3) v);
    method Action S_AXI_HP3_ARVALID(Bit#(1) v);
    method Action S_AXI_HP3_AWADDR(Bit#(32) v);
    method Action S_AXI_HP3_AWBURST(Bit#(2) v);
    method Action S_AXI_HP3_AWCACHE(Bit#(4) v);
    method Action S_AXI_HP3_AWID(Bit#(C_S_AXI_HP3_ID_WIDTH) v);
    method Action S_AXI_HP3_AWLEN(Bit#(4) v);
    method Action S_AXI_HP3_AWLOCK(Bit#(2) v);
    method Action S_AXI_HP3_AWPROT(Bit#(3) v);
    method Action S_AXI_HP3_AWQOS(Bit#(4) v);
    method Bit#(1) S_AXI_HP3_AWREADY();
    method Action S_AXI_HP3_AWSIZE(Bit#(3) v);
    method Action S_AXI_HP3_AWVALID(Bit#(1) v);
    method Bit#(C_S_AXI_HP3_ID_WIDTH) S_AXI_HP3_BID();
    method Action S_AXI_HP3_BREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP3_BRESP();
    method Bit#(1) S_AXI_HP3_BVALID();
    method Bit#(3) S_AXI_HP3_RACOUNT();
    method Bit#(8) S_AXI_HP3_RCOUNT();
    method Bit#(C_S_AXI_HP3_DATA_WIDTH) S_AXI_HP3_RDATA();
    method Action S_AXI_HP3_RDISSUECAP1_EN(Bit#(1) v);
    method Bit#(C_S_AXI_HP3_ID_WIDTH) S_AXI_HP3_RID();
    method Bit#(1) S_AXI_HP3_RLAST();
    method Action S_AXI_HP3_RREADY(Bit#(1) v);
    method Bit#(2) S_AXI_HP3_RRESP();
    method Bit#(1) S_AXI_HP3_RVALID();
    method Bit#(6) S_AXI_HP3_WACOUNT();
    method Bit#(8) S_AXI_HP3_WCOUNT();
    method Action S_AXI_HP3_WDATA(Bit#(C_S_AXI_HP3_DATA_WIDTH) v);
    method Action S_AXI_HP3_WID(Bit#(C_S_AXI_HP3_ID_WIDTH) v);
    method Action S_AXI_HP3_WLAST(Bit#(1) v);
    method Bit#(1) S_AXI_HP3_WREADY();
    method Action S_AXI_HP3_WRISSUECAP1_EN(Bit#(1) v);
    method Action S_AXI_HP3_WSTRB(Bit#(C_S_AXI_HP3_DATA_WIDTH/8) v);
    method Action S_AXI_HP3_WVALID(Bit#(1) v);
    method Action TRACE_CLK(Bit#(1) v);
    method Bit#(1) TRACE_CTL();
    method Bit#(32) TRACE_DATA();
    method Action TTC0_CLK0_IN(Bit#(1) v);
    method Action TTC0_CLK1_IN(Bit#(1) v);
    method Action TTC0_CLK2_IN(Bit#(1) v);
    method Bit#(1) TTC0_WAVE0_OUT();
    method Bit#(1) TTC0_WAVE1_OUT();
    method Bit#(1) TTC0_WAVE2_OUT();
    method Action TTC1_CLK0_IN(Bit#(1) v);
    method Action TTC1_CLK1_IN(Bit#(1) v);
    method Action TTC1_CLK2_IN(Bit#(1) v);
    method Bit#(1) TTC1_WAVE0_OUT();
    method Bit#(1) TTC1_WAVE1_OUT();
    method Bit#(1) TTC1_WAVE2_OUT();
    method Action UART0_CTSN(Bit#(1) v);
    method Action UART0_DCDN(Bit#(1) v);
    method Action UART0_DSRN(Bit#(1) v);
    method Bit#(1) UART0_DTRN();
    method Action UART0_RIN(Bit#(1) v);
    method Bit#(1) UART0_RTSN();
    method Action UART0_RX(Bit#(1) v);
    method Bit#(1) UART0_TX();
    method Action UART1_CTSN(Bit#(1) v);
    method Action UART1_DCDN(Bit#(1) v);
    method Action UART1_DSRN(Bit#(1) v);
    method Bit#(1) UART1_DTRN();
    method Action UART1_RIN(Bit#(1) v);
    method Bit#(1) UART1_RTSN();
    method Action UART1_RX(Bit#(1) v);
    method Bit#(1) UART1_TX();
    method Bit#(2) USB0_PORT_INDCTL();
    method Action USB0_VBUS_PWRFAULT(Bit#(1) v);
    method Bit#(1) USB0_VBUS_PWRSELECT();
    method Bit#(2) USB1_PORT_INDCTL();
    method Action USB1_VBUS_PWRFAULT(Bit#(1) v);
    method Bit#(1) USB1_VBUS_PWRSELECT();
    method Action WDT_CLK_IN(Bit#(1) v);
    method Bit#(1) WDT_RST_OUT();

   schedule (datain, idatain, inc, ce) CF (datain, idatain, inc, ce);
endmodule
