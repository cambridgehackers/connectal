//Top.bsv customized for Ring example

// bsv libraries
import Vector::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import Portal::*;
import AxiMasterSlave::*;
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;


// generated by tool
import RingIndicationProxy::*;
import RingRequestWrapper::*;

// defined by user
import Ring::*;

module mkPortalTop(StdPortalTop);

   // instantiate user portals
   RingIndicationProxy echoIndicationProxy <- mkRingIndicationProxy(7);
   RingRequestInternal echoRequestInternal <- mkRingRequestInternal(echoIndicationProxy.ifc);
   RingRequestWrapper echoRequestWrapper <- mkRingRequestWrapper(1008,echoRequestInternal.ifc);
   
   
   Vector#(2,StdPortal) portals;
   portals[0] = echoIndicationProxy.portalIfc;
   portals[1] = echoRequestWrapper.portalIfc; 

   let interrupt_mux <- mkInterruptMux(portals);
   
   // instantiate system directory
   Directory dir <- mkDirectoryDbg(portals,interrupt_mux);
   Vector#(1,StdPortal) directories;
   directories[0] = dir.portalIfc;
   
   // when constructing the ctrl mux, directories must be the first argument
   let ctrl_mux <- mkAxiSlaveMux(directories,portals);
   
   interface ReadOnly interrupt = interrupt_mux;
   interface StdAxi3Slave ctrl = ctrl_mux;


endmodule : mkPortalTop
