
// Copyright (c) 2013 Nokia, Inc.
// Copyright (c) 2013 Quanta Research Cambridge, Inc.

// Permission is hereby granted, free of charge, to any person
// obtaining a copy of this software and associated documentation
// files (the "Software"), to deal in the Software without
// restriction, including without limitation the rights to use, copy,
// modify, merge, publish, distribute, sublicense, and/or sell copies
// of the Software, and to permit persons to whom the Software is
// furnished to do so, subject to the following conditions:

// The above copyright notice and this permission notice shall be
// included in all copies or substantial portions of the Software.

// THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND,
// EXPRESS OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF
// MERCHANTABILITY, FITNESS FOR A PARTICULAR PURPOSE AND
// NONINFRINGEMENT. IN NO EVENT SHALL THE AUTHORS OR COPYRIGHT HOLDERS
// BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER LIABILITY, WHETHER IN AN
// ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING FROM, OUT OF OR IN
// CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER DEALINGS IN THE
// SOFTWARE.

import Vector            :: *;
import Clocks            :: *;
import Connectable       :: *;
import Assert            :: *;
import Xilinx            :: *;
import XilinxPCIE        :: *;
import Xilinx7PcieBridge :: *;
import PcieToAxiBridge   :: *;

import Echo::*;

// the following three are generated by the script from the interface declarations
import CoreEchoRequestWrapper::*;
import NonEchoRequestWrapper::*;
import CoreEchoIndicationProxy::*;

import AxiMasterSlave::*;
import AxiClientServer::*;

module mkEchoPcie#(X7PcieBridgeIfc#(8) x7pcie)(KC705_FPGA);

   CoreEchoIndicationProxy coreIndicationProxy <- mkCoreEchoIndicationProxy();

   EchoRequest echoRequest <- mkEchoRequest( coreIndicationProxy );

   CoreEchoRequestWrapper coreRequestWrapper <- mkCoreEchoRequestWrapper(echoRequest.coreRequest);
   NonEchoRequestWrapper otherRequestWrapper <- mkNonEchoRequestWrapper(echoRequest.otherRequest);

   Vector#(numPortals,Axi3Slave#(32,32,4,12)) ctrls_v;
   ctrls_v[0] = coreIndicationProxy.ctrl;
   ctrls_v[1] = coreRequestWrapper.ctrl;
   ctrls_v[2] = coreRequestWrapper.ctrl;
   let ctrl_mux <- mkAxiSlaveMux(ctrls_v);
   mkConnection(x7pcie.portal0, ctrl_mux);

   Vector#(numPortals,ReadOnly#(Bool)) interrupts_v;
   interrupts_v[0] = coreIndicationProxy.interrupt;
   interrupts_v[1] = coreRequestWrapper.interrupt;
   interrupts_v[2] = otherRequestWrapper.interrupt;
   mkConnection(x7pcie.interrupts, interrupts_v);

   interface pcie = x7pcie.pcie;
   method leds = zeroExtend({  pack(x7pcie.isCalibrated)
			     , pack(True)
			     , pack(False)
			     , pack(x7pcie.isLinkUp)
			     });
endmodule

(* synthesize, no_default_clock, no_default_reset *)
module mkEchoPcieTop #(Clock pci_sys_clk_p, Clock pci_sys_clk_n,
                          Clock sys_clk_p,     Clock sys_clk_n,
                          Reset pci_sys_reset_n)
                         (KC705_FPGA);

   let contentId = 64'h4563686f;
   let numPortals = 3;
   X7PcieBridgeIfc#(8) x7pcie <- mkX7PcieBridge(pci_sys_clk_p, pci_sys_clk_n, sys_clk_p, sys_clk_n, pci_sys_reset_n,
						numPortals,
						contentId );

   let top <- mkEchoPcie(x7pcie, clocked_by x7pcie.clock125, reset_by x7pcie.reset125);
   interface pcie = top.pcie;
   methods leds = top.leds;
   
endmodule: mkEchoPcieTop
