import Clocks::*;
import DefaultValue::*;

import "BVI" test_program =
module mkTestProgram(Empty);
    default_clock clk();
    default_reset rst();
endmodule
