// bsv libraries
import SpecialFIFOs::*;
import Vector::*;
import StmtFSM::*;
import FIFO::*;
import Connectable::*;

// portz libraries
import Directory::*;
import CtrlMux::*;
import Portal::*;
import Leds::*;
import PortalMemory::*;
import MemServer::*;
import SGList::*;
import PortalMemory::*;
import MemTypes::*;
import MemUtils::*;
import RbmTypes::*;
import HostInterface::*;

// generated by tool
import DmaDebugRequestWrapper::*;
import SGListConfigRequestWrapper::*;
import DmaDebugIndicationProxy::*;
import SGListConfigIndicationProxy::*;

module  mkPortalTop#(HostType host)(PortalTop#(PhysAddrWidth,TMul#(32,N),Empty,NumberOfMasters));

   // all this stuff is here so we can call portalAlloc in user space
   let reader <- mkMemReader();
   let writer <- mkMemWriter();

   Vector#(1,ObjectReadClient#(TMul#(32,N)))  readClients  = cons(reader.readClient, nil);
   Vector#(1,ObjectWriteClient#(TMul#(32,N))) writeClients = cons(writer.writeClient, nil);

   SGListConfigIndicationProxy hostmemSGListConfigIndicationProxy <- mkSGListConfigIndicationProxy(HostmemSGListConfigIndication);
   SGListMMU#(PhysAddrWidth) hostmemSGList <- mkSGListMMU(0, True, hostmemSGListConfigIndicationProxy.ifc);
   SGListConfigRequestWrapper hostmemSGListConfigRequestWrapper <- mkSGListConfigRequestWrapper(HostmemSGListConfigRequest, hostmemSGList.request);

   DmaDebugIndicationProxy hostmemDmaDebugIndicationProxy <- mkDmaDebugIndicationProxy(HostmemDmaDebugIndication);
   MemServer#(PhysAddrWidth,TMul#(32,N), NumberOfMasters) dma <- mkMemServerRW(hostmemDmaDebugIndicationProxy.ifc, readClients, writeClients, cons(hostmemSGList,nil));
   DmaDebugRequestWrapper hostmemDmaDebugRequestWrapper <- mkDmaDebugRequestWrapper(HostmemDmaDebugRequest, dma.request);

   Vector#(4,StdPortal) portals;
   portals[0] = hostmemDmaDebugIndicationProxy.portalIfc; 
   portals[1] = hostmemDmaDebugRequestWrapper.portalIfc;
   portals[2] = hostmemSGListConfigRequestWrapper.portalIfc;
   portals[3] = hostmemSGListConfigIndicationProxy.portalIfc;


   StdDirectory dir <- mkStdDirectory(portals);
   let ctrl_mux <- mkSlaveMux(dir,portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;

endmodule : mkPortalTop
