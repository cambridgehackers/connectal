/* Copyright (c) 2014 Quanta Research Cambridge, Inc
 *
 * Permission is hereby granted, free of charge, to any person obtaining a
 * copy of this software and associated documentation files (the "Software"),
 * to deal in the Software without restriction, including without limitation
 * the rights to use, copy, modify, merge, publish, distribute, sublicense,
 * and/or sell copies of the Software, and to permit persons to whom the
 * Software is furnished to do so, subject to the following conditions:
 *
 * The above copyright notice and this permission notice shall be included
 * in all copies or substantial portions of the Software.
 *
 * THE SOFTWARE IS PROVIDED "AS IS", WITHOUT WARRANTY OF ANY KIND, EXPRESS
 * OR IMPLIED, INCLUDING BUT NOT LIMITED TO THE WARRANTIES OF MERCHANTABILITY,
 * FITNESS FOR A PARTICULAR PURPOSE AND NONINFRINGEMENT. IN NO EVENT SHALL
 * THE AUTHORS OR COPYRIGHT HOLDERS BE LIABLE FOR ANY CLAIM, DAMAGES OR OTHER
 * LIABILITY, WHETHER IN AN ACTION OF CONTRACT, TORT OR OTHERWISE, ARISING
 * FROM, OUT OF OR IN CONNECTION WITH THE SOFTWARE OR THE USE OR OTHER
 * DEALINGS IN THE SOFTWARE.
 */
import Vector::*;
import FIFO::*;
import Connectable::*;
import CtrlMux::*;
import Portal::*;
import HostInterface::*;
import Leds::*;
import MMU::*;
import MemServer::*;
import MemPortal::*;
import SharedMemoryPortal::*;

// generated by tool
import Simple::*;
import SimpleRequest::*;
import MMURequest::*;
import MMUIndication::*;
import SharedMemoryPortalConfig::*;
import MemServerIndication::*;

// defined by user
import Simple::*;

typedef enum {SimpleRequestH2S, SimpleRequestS2H,
	      MMURequestS2H, MMUIndicationH2S, MemServerIndicationH2S, ReqConfigWrapper, IndConfigWrapper} IfcNames deriving (Eq,Bits);

module mkConnectalTop(StdConnectalDmaTop#(PhysAddrWidth));

   // instantiate DUT
   SimpleRequestProxyPortal lSimpleRequestProxyPortal <- mkSimpleRequestProxyPortal(SimpleRequestH2S);
   SharedMemoryPortal#(64) lSimpleRequestProxyPortalMem <- mkSharedMemoryPortal(lSimpleRequestProxyPortal.portalIfc);
   SharedMemoryPortalConfigWrapper lSimpleRequestProxy <-
       mkSharedMemoryPortalConfigWrapper(IndConfigWrapper, lSimpleRequestProxyPortalMem.cfg);
   //SimpleRequestProxy lSimpleRequestProxy <- mkSimpleRequestProxy(SimpleRequestH2S);

   Simple lSimple <- mkSimple(lSimpleRequestProxyPortal.ifc);
   //Simple lSimple <- mkSimple(lSimpleRequestProxy.ifc);

   SimpleRequestWrapperPortal lSimpleRequestWrapperPortal <- mkSimpleRequestWrapperPortal(SimpleRequestS2H,lSimple.request);
   SharedMemoryPortal#(64) lSimpleRequestWrapperPortalMem <- mkSharedMemoryPortal(lSimpleRequestWrapperPortal.portalIfc);
   SharedMemoryPortalConfigWrapper lSimpleRequestWrapper <-
       mkSharedMemoryPortalConfigWrapper(ReqConfigWrapper, lSimpleRequestWrapperPortalMem.cfg);
   //SimpleRequestWrapper lSimpleRequestWrapper <- mkSimpleRequestWrapper(SimpleRequestS2H, lSimple.request);

   // MMU used for shared memory buffer mapping
   MMUIndicationProxy lMMUIndicationProxy <- mkMMUIndicationProxy(MMUIndicationH2S);
   MMU#(PhysAddrWidth) mmu <- mkMMU(0, True, lMMUIndicationProxy.ifc);
   MMURequestWrapper lMMURequestWrapper <- mkMMURequestWrapper(MMURequestS2H, mmu.request);

   // MemServer used for shared memory buffer access
   MemServerIndicationProxy lMemServerIndicationProxy <- mkMemServerIndicationProxy(MemServerIndicationH2S);
   MemServer#(PhysAddrWidth,64,1) dma <- mkMemServerRW(lMemServerIndicationProxy.ifc,
       cons(lSimpleRequestWrapperPortalMem.readClient,cons(lSimpleRequestProxyPortalMem.readClient,nil)),
       cons(lSimpleRequestWrapperPortalMem.writeClient,cons(lSimpleRequestProxyPortalMem.writeClient,nil)), cons(mmu,nil));

   Vector#(5,StdPortal) portals;
   portals[0] = lMMURequestWrapper.portalIfc;
   portals[1] = lMMUIndicationProxy.portalIfc;
   portals[2] = lSimpleRequestWrapper.portalIfc;
   portals[3] = lSimpleRequestProxy.portalIfc;
   portals[4] = lMemServerIndicationProxy.portalIfc;
   let ctrl_mux <- mkSlaveMux(portals);
   
   interface interrupt = getInterruptVector(portals);
   interface slave = ctrl_mux;
   interface masters = dma.masters;
   interface leds = default_leds;
endmodule : mkConnectalTop
