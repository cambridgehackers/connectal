
typeclass PortalMemory#(type a);
endtypeclass
   